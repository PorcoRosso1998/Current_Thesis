module Tables();
	reg [13:0] logarithm_table[8191:0];
	reg [13:0] Dplus[8191:0];
	reg [13:0] Dminus[8191:0];
	initial begin
		logarithm_table[1] = 14'b1111001_0000000;
		logarithm_table[2] = 14'b1111010_0000000;
		logarithm_table[3] = 14'b1111010_1001011;
		logarithm_table[4] = 14'b1111011_0000000;
		logarithm_table[5] = 14'b1111011_0101001;
		logarithm_table[6] = 14'b1111011_1001011;
		logarithm_table[7] = 14'b1111011_1100111;
		logarithm_table[8] = 14'b1111100_0000000;
		logarithm_table[9] = 14'b1111100_0010110;
		logarithm_table[10] = 14'b1111100_0101001;
		logarithm_table[11] = 14'b1111100_0111011;
		logarithm_table[12] = 14'b1111100_1001011;
		logarithm_table[13] = 14'b1111100_1011010;
		logarithm_table[14] = 14'b1111100_1100111;
		logarithm_table[15] = 14'b1111100_1110100;
		logarithm_table[16] = 14'b1111101_0000000;
		logarithm_table[17] = 14'b1111101_0001011;
		logarithm_table[18] = 14'b1111101_0010110;
		logarithm_table[19] = 14'b1111101_0100000;
		logarithm_table[20] = 14'b1111101_0101001;
		logarithm_table[21] = 14'b1111101_0110010;
		logarithm_table[22] = 14'b1111101_0111011;
		logarithm_table[23] = 14'b1111101_1000011;
		logarithm_table[24] = 14'b1111101_1001011;
		logarithm_table[25] = 14'b1111101_1010010;
		logarithm_table[26] = 14'b1111101_1011010;
		logarithm_table[27] = 14'b1111101_1100001;
		logarithm_table[28] = 14'b1111101_1100111;
		logarithm_table[29] = 14'b1111101_1101110;
		logarithm_table[30] = 14'b1111101_1110100;
		logarithm_table[31] = 14'b1111101_1111010;
		logarithm_table[32] = 14'b1111110_0000000;
		logarithm_table[33] = 14'b1111110_0000110;
		logarithm_table[34] = 14'b1111110_0001011;
		logarithm_table[35] = 14'b1111110_0010001;
		logarithm_table[36] = 14'b1111110_0010110;
		logarithm_table[37] = 14'b1111110_0011011;
		logarithm_table[38] = 14'b1111110_0100000;
		logarithm_table[39] = 14'b1111110_0100101;
		logarithm_table[40] = 14'b1111110_0101001;
		logarithm_table[41] = 14'b1111110_0101110;
		logarithm_table[42] = 14'b1111110_0110010;
		logarithm_table[43] = 14'b1111110_0110111;
		logarithm_table[44] = 14'b1111110_0111011;
		logarithm_table[45] = 14'b1111110_0111111;
		logarithm_table[46] = 14'b1111110_1000011;
		logarithm_table[47] = 14'b1111110_1000111;
		logarithm_table[48] = 14'b1111110_1001011;
		logarithm_table[49] = 14'b1111110_1001111;
		logarithm_table[50] = 14'b1111110_1010010;
		logarithm_table[51] = 14'b1111110_1010110;
		logarithm_table[52] = 14'b1111110_1011010;
		logarithm_table[53] = 14'b1111110_1011101;
		logarithm_table[54] = 14'b1111110_1100001;
		logarithm_table[55] = 14'b1111110_1100100;
		logarithm_table[56] = 14'b1111110_1100111;
		logarithm_table[57] = 14'b1111110_1101011;
		logarithm_table[58] = 14'b1111110_1101110;
		logarithm_table[59] = 14'b1111110_1110001;
		logarithm_table[60] = 14'b1111110_1110100;
		logarithm_table[61] = 14'b1111110_1110111;
		logarithm_table[62] = 14'b1111110_1111010;
		logarithm_table[63] = 14'b1111110_1111101;
		logarithm_table[64] = 14'b1111111_0000000;
		logarithm_table[65] = 14'b1111111_0000011;
		logarithm_table[66] = 14'b1111111_0000110;
		logarithm_table[67] = 14'b1111111_0001000;
		logarithm_table[68] = 14'b1111111_0001011;
		logarithm_table[69] = 14'b1111111_0001110;
		logarithm_table[70] = 14'b1111111_0010001;
		logarithm_table[71] = 14'b1111111_0010011;
		logarithm_table[72] = 14'b1111111_0010110;
		logarithm_table[73] = 14'b1111111_0011000;
		logarithm_table[74] = 14'b1111111_0011011;
		logarithm_table[75] = 14'b1111111_0011101;
		logarithm_table[76] = 14'b1111111_0100000;
		logarithm_table[77] = 14'b1111111_0100010;
		logarithm_table[78] = 14'b1111111_0100101;
		logarithm_table[79] = 14'b1111111_0100111;
		logarithm_table[80] = 14'b1111111_0101001;
		logarithm_table[81] = 14'b1111111_0101100;
		logarithm_table[82] = 14'b1111111_0101110;
		logarithm_table[83] = 14'b1111111_0110000;
		logarithm_table[84] = 14'b1111111_0110010;
		logarithm_table[85] = 14'b1111111_0110100;
		logarithm_table[86] = 14'b1111111_0110111;
		logarithm_table[87] = 14'b1111111_0111001;
		logarithm_table[88] = 14'b1111111_0111011;
		logarithm_table[89] = 14'b1111111_0111101;
		logarithm_table[90] = 14'b1111111_0111111;
		logarithm_table[91] = 14'b1111111_1000001;
		logarithm_table[92] = 14'b1111111_1000011;
		logarithm_table[93] = 14'b1111111_1000101;
		logarithm_table[94] = 14'b1111111_1000111;
		logarithm_table[95] = 14'b1111111_1001001;
		logarithm_table[96] = 14'b1111111_1001011;
		logarithm_table[97] = 14'b1111111_1001101;
		logarithm_table[98] = 14'b1111111_1001111;
		logarithm_table[99] = 14'b1111111_1010001;
		logarithm_table[100] = 14'b1111111_1010010;
		logarithm_table[101] = 14'b1111111_1010100;
		logarithm_table[102] = 14'b1111111_1010110;
		logarithm_table[103] = 14'b1111111_1011000;
		logarithm_table[104] = 14'b1111111_1011010;
		logarithm_table[105] = 14'b1111111_1011011;
		logarithm_table[106] = 14'b1111111_1011101;
		logarithm_table[107] = 14'b1111111_1011111;
		logarithm_table[108] = 14'b1111111_1100001;
		logarithm_table[109] = 14'b1111111_1100010;
		logarithm_table[110] = 14'b1111111_1100100;
		logarithm_table[111] = 14'b1111111_1100110;
		logarithm_table[112] = 14'b1111111_1100111;
		logarithm_table[113] = 14'b1111111_1101001;
		logarithm_table[114] = 14'b1111111_1101011;
		logarithm_table[115] = 14'b1111111_1101100;
		logarithm_table[116] = 14'b1111111_1101110;
		logarithm_table[117] = 14'b1111111_1101111;
		logarithm_table[118] = 14'b1111111_1110001;
		logarithm_table[119] = 14'b1111111_1110011;
		logarithm_table[120] = 14'b1111111_1110100;
		logarithm_table[121] = 14'b1111111_1110110;
		logarithm_table[122] = 14'b1111111_1110111;
		logarithm_table[123] = 14'b1111111_1111001;
		logarithm_table[124] = 14'b1111111_1111010;
		logarithm_table[125] = 14'b1111111_1111100;
		logarithm_table[126] = 14'b1111111_1111101;
		logarithm_table[127] = 14'b1111111_1111111;
		logarithm_table[128] = 14'b0000000_0000000;
		logarithm_table[129] = 14'b0000000_0000001;
		logarithm_table[130] = 14'b0000000_0000011;
		logarithm_table[131] = 14'b0000000_0000100;
		logarithm_table[132] = 14'b0000000_0000110;
		logarithm_table[133] = 14'b0000000_0000111;
		logarithm_table[134] = 14'b0000000_0001000;
		logarithm_table[135] = 14'b0000000_0001010;
		logarithm_table[136] = 14'b0000000_0001011;
		logarithm_table[137] = 14'b0000000_0001101;
		logarithm_table[138] = 14'b0000000_0001110;
		logarithm_table[139] = 14'b0000000_0001111;
		logarithm_table[140] = 14'b0000000_0010001;
		logarithm_table[141] = 14'b0000000_0010010;
		logarithm_table[142] = 14'b0000000_0010011;
		logarithm_table[143] = 14'b0000000_0010100;
		logarithm_table[144] = 14'b0000000_0010110;
		logarithm_table[145] = 14'b0000000_0010111;
		logarithm_table[146] = 14'b0000000_0011000;
		logarithm_table[147] = 14'b0000000_0011010;
		logarithm_table[148] = 14'b0000000_0011011;
		logarithm_table[149] = 14'b0000000_0011100;
		logarithm_table[150] = 14'b0000000_0011101;
		logarithm_table[151] = 14'b0000000_0011111;
		logarithm_table[152] = 14'b0000000_0100000;
		logarithm_table[153] = 14'b0000000_0100001;
		logarithm_table[154] = 14'b0000000_0100010;
		logarithm_table[155] = 14'b0000000_0100011;
		logarithm_table[156] = 14'b0000000_0100101;
		logarithm_table[157] = 14'b0000000_0100110;
		logarithm_table[158] = 14'b0000000_0100111;
		logarithm_table[159] = 14'b0000000_0101000;
		logarithm_table[160] = 14'b0000000_0101001;
		logarithm_table[161] = 14'b0000000_0101010;
		logarithm_table[162] = 14'b0000000_0101100;
		logarithm_table[163] = 14'b0000000_0101101;
		logarithm_table[164] = 14'b0000000_0101110;
		logarithm_table[165] = 14'b0000000_0101111;
		logarithm_table[166] = 14'b0000000_0110000;
		logarithm_table[167] = 14'b0000000_0110001;
		logarithm_table[168] = 14'b0000000_0110010;
		logarithm_table[169] = 14'b0000000_0110011;
		logarithm_table[170] = 14'b0000000_0110100;
		logarithm_table[171] = 14'b0000000_0110101;
		logarithm_table[172] = 14'b0000000_0110111;
		logarithm_table[173] = 14'b0000000_0111000;
		logarithm_table[174] = 14'b0000000_0111001;
		logarithm_table[175] = 14'b0000000_0111010;
		logarithm_table[176] = 14'b0000000_0111011;
		logarithm_table[177] = 14'b0000000_0111100;
		logarithm_table[178] = 14'b0000000_0111101;
		logarithm_table[179] = 14'b0000000_0111110;
		logarithm_table[180] = 14'b0000000_0111111;
		logarithm_table[181] = 14'b0000000_1000000;
		logarithm_table[182] = 14'b0000000_1000001;
		logarithm_table[183] = 14'b0000000_1000010;
		logarithm_table[184] = 14'b0000000_1000011;
		logarithm_table[185] = 14'b0000000_1000100;
		logarithm_table[186] = 14'b0000000_1000101;
		logarithm_table[187] = 14'b0000000_1000110;
		logarithm_table[188] = 14'b0000000_1000111;
		logarithm_table[189] = 14'b0000000_1001000;
		logarithm_table[190] = 14'b0000000_1001001;
		logarithm_table[191] = 14'b0000000_1001010;
		logarithm_table[192] = 14'b0000000_1001011;
		logarithm_table[193] = 14'b0000000_1001100;
		logarithm_table[194] = 14'b0000000_1001101;
		logarithm_table[195] = 14'b0000000_1001110;
		logarithm_table[196] = 14'b0000000_1001111;
		logarithm_table[197] = 14'b0000000_1010000;
		logarithm_table[198] = 14'b0000000_1010001;
		logarithm_table[199] = 14'b0000000_1010001;
		logarithm_table[200] = 14'b0000000_1010010;
		logarithm_table[201] = 14'b0000000_1010011;
		logarithm_table[202] = 14'b0000000_1010100;
		logarithm_table[203] = 14'b0000000_1010101;
		logarithm_table[204] = 14'b0000000_1010110;
		logarithm_table[205] = 14'b0000000_1010111;
		logarithm_table[206] = 14'b0000000_1011000;
		logarithm_table[207] = 14'b0000000_1011001;
		logarithm_table[208] = 14'b0000000_1011010;
		logarithm_table[209] = 14'b0000000_1011011;
		logarithm_table[210] = 14'b0000000_1011011;
		logarithm_table[211] = 14'b0000000_1011100;
		logarithm_table[212] = 14'b0000000_1011101;
		logarithm_table[213] = 14'b0000000_1011110;
		logarithm_table[214] = 14'b0000000_1011111;
		logarithm_table[215] = 14'b0000000_1100000;
		logarithm_table[216] = 14'b0000000_1100001;
		logarithm_table[217] = 14'b0000000_1100001;
		logarithm_table[218] = 14'b0000000_1100010;
		logarithm_table[219] = 14'b0000000_1100011;
		logarithm_table[220] = 14'b0000000_1100100;
		logarithm_table[221] = 14'b0000000_1100101;
		logarithm_table[222] = 14'b0000000_1100110;
		logarithm_table[223] = 14'b0000000_1100111;
		logarithm_table[224] = 14'b0000000_1100111;
		logarithm_table[225] = 14'b0000000_1101000;
		logarithm_table[226] = 14'b0000000_1101001;
		logarithm_table[227] = 14'b0000000_1101010;
		logarithm_table[228] = 14'b0000000_1101011;
		logarithm_table[229] = 14'b0000000_1101011;
		logarithm_table[230] = 14'b0000000_1101100;
		logarithm_table[231] = 14'b0000000_1101101;
		logarithm_table[232] = 14'b0000000_1101110;
		logarithm_table[233] = 14'b0000000_1101111;
		logarithm_table[234] = 14'b0000000_1101111;
		logarithm_table[235] = 14'b0000000_1110000;
		logarithm_table[236] = 14'b0000000_1110001;
		logarithm_table[237] = 14'b0000000_1110010;
		logarithm_table[238] = 14'b0000000_1110011;
		logarithm_table[239] = 14'b0000000_1110011;
		logarithm_table[240] = 14'b0000000_1110100;
		logarithm_table[241] = 14'b0000000_1110101;
		logarithm_table[242] = 14'b0000000_1110110;
		logarithm_table[243] = 14'b0000000_1110110;
		logarithm_table[244] = 14'b0000000_1110111;
		logarithm_table[245] = 14'b0000000_1111000;
		logarithm_table[246] = 14'b0000000_1111001;
		logarithm_table[247] = 14'b0000000_1111001;
		logarithm_table[248] = 14'b0000000_1111010;
		logarithm_table[249] = 14'b0000000_1111011;
		logarithm_table[250] = 14'b0000000_1111100;
		logarithm_table[251] = 14'b0000000_1111100;
		logarithm_table[252] = 14'b0000000_1111101;
		logarithm_table[253] = 14'b0000000_1111110;
		logarithm_table[254] = 14'b0000000_1111111;
		logarithm_table[255] = 14'b0000000_1111111;
		logarithm_table[256] = 14'b0000001_0000000;
		logarithm_table[257] = 14'b0000001_0000001;
		logarithm_table[258] = 14'b0000001_0000001;
		logarithm_table[259] = 14'b0000001_0000010;
		logarithm_table[260] = 14'b0000001_0000011;
		logarithm_table[261] = 14'b0000001_0000100;
		logarithm_table[262] = 14'b0000001_0000100;
		logarithm_table[263] = 14'b0000001_0000101;
		logarithm_table[264] = 14'b0000001_0000110;
		logarithm_table[265] = 14'b0000001_0000110;
		logarithm_table[266] = 14'b0000001_0000111;
		logarithm_table[267] = 14'b0000001_0001000;
		logarithm_table[268] = 14'b0000001_0001000;
		logarithm_table[269] = 14'b0000001_0001001;
		logarithm_table[270] = 14'b0000001_0001010;
		logarithm_table[271] = 14'b0000001_0001011;
		logarithm_table[272] = 14'b0000001_0001011;
		logarithm_table[273] = 14'b0000001_0001100;
		logarithm_table[274] = 14'b0000001_0001101;
		logarithm_table[275] = 14'b0000001_0001101;
		logarithm_table[276] = 14'b0000001_0001110;
		logarithm_table[277] = 14'b0000001_0001111;
		logarithm_table[278] = 14'b0000001_0001111;
		logarithm_table[279] = 14'b0000001_0010000;
		logarithm_table[280] = 14'b0000001_0010001;
		logarithm_table[281] = 14'b0000001_0010001;
		logarithm_table[282] = 14'b0000001_0010010;
		logarithm_table[283] = 14'b0000001_0010011;
		logarithm_table[284] = 14'b0000001_0010011;
		logarithm_table[285] = 14'b0000001_0010100;
		logarithm_table[286] = 14'b0000001_0010100;
		logarithm_table[287] = 14'b0000001_0010101;
		logarithm_table[288] = 14'b0000001_0010110;
		logarithm_table[289] = 14'b0000001_0010110;
		logarithm_table[290] = 14'b0000001_0010111;
		logarithm_table[291] = 14'b0000001_0011000;
		logarithm_table[292] = 14'b0000001_0011000;
		logarithm_table[293] = 14'b0000001_0011001;
		logarithm_table[294] = 14'b0000001_0011010;
		logarithm_table[295] = 14'b0000001_0011010;
		logarithm_table[296] = 14'b0000001_0011011;
		logarithm_table[297] = 14'b0000001_0011011;
		logarithm_table[298] = 14'b0000001_0011100;
		logarithm_table[299] = 14'b0000001_0011101;
		logarithm_table[300] = 14'b0000001_0011101;
		logarithm_table[301] = 14'b0000001_0011110;
		logarithm_table[302] = 14'b0000001_0011111;
		logarithm_table[303] = 14'b0000001_0011111;
		logarithm_table[304] = 14'b0000001_0100000;
		logarithm_table[305] = 14'b0000001_0100000;
		logarithm_table[306] = 14'b0000001_0100001;
		logarithm_table[307] = 14'b0000001_0100010;
		logarithm_table[308] = 14'b0000001_0100010;
		logarithm_table[309] = 14'b0000001_0100011;
		logarithm_table[310] = 14'b0000001_0100011;
		logarithm_table[311] = 14'b0000001_0100100;
		logarithm_table[312] = 14'b0000001_0100101;
		logarithm_table[313] = 14'b0000001_0100101;
		logarithm_table[314] = 14'b0000001_0100110;
		logarithm_table[315] = 14'b0000001_0100110;
		logarithm_table[316] = 14'b0000001_0100111;
		logarithm_table[317] = 14'b0000001_0100111;
		logarithm_table[318] = 14'b0000001_0101000;
		logarithm_table[319] = 14'b0000001_0101001;
		logarithm_table[320] = 14'b0000001_0101001;
		logarithm_table[321] = 14'b0000001_0101010;
		logarithm_table[322] = 14'b0000001_0101010;
		logarithm_table[323] = 14'b0000001_0101011;
		logarithm_table[324] = 14'b0000001_0101100;
		logarithm_table[325] = 14'b0000001_0101100;
		logarithm_table[326] = 14'b0000001_0101101;
		logarithm_table[327] = 14'b0000001_0101101;
		logarithm_table[328] = 14'b0000001_0101110;
		logarithm_table[329] = 14'b0000001_0101110;
		logarithm_table[330] = 14'b0000001_0101111;
		logarithm_table[331] = 14'b0000001_0101111;
		logarithm_table[332] = 14'b0000001_0110000;
		logarithm_table[333] = 14'b0000001_0110001;
		logarithm_table[334] = 14'b0000001_0110001;
		logarithm_table[335] = 14'b0000001_0110010;
		logarithm_table[336] = 14'b0000001_0110010;
		logarithm_table[337] = 14'b0000001_0110011;
		logarithm_table[338] = 14'b0000001_0110011;
		logarithm_table[339] = 14'b0000001_0110100;
		logarithm_table[340] = 14'b0000001_0110100;
		logarithm_table[341] = 14'b0000001_0110101;
		logarithm_table[342] = 14'b0000001_0110101;
		logarithm_table[343] = 14'b0000001_0110110;
		logarithm_table[344] = 14'b0000001_0110111;
		logarithm_table[345] = 14'b0000001_0110111;
		logarithm_table[346] = 14'b0000001_0111000;
		logarithm_table[347] = 14'b0000001_0111000;
		logarithm_table[348] = 14'b0000001_0111001;
		logarithm_table[349] = 14'b0000001_0111001;
		logarithm_table[350] = 14'b0000001_0111010;
		logarithm_table[351] = 14'b0000001_0111010;
		logarithm_table[352] = 14'b0000001_0111011;
		logarithm_table[353] = 14'b0000001_0111011;
		logarithm_table[354] = 14'b0000001_0111100;
		logarithm_table[355] = 14'b0000001_0111100;
		logarithm_table[356] = 14'b0000001_0111101;
		logarithm_table[357] = 14'b0000001_0111101;
		logarithm_table[358] = 14'b0000001_0111110;
		logarithm_table[359] = 14'b0000001_0111110;
		logarithm_table[360] = 14'b0000001_0111111;
		logarithm_table[361] = 14'b0000001_0111111;
		logarithm_table[362] = 14'b0000001_1000000;
		logarithm_table[363] = 14'b0000001_1000000;
		logarithm_table[364] = 14'b0000001_1000001;
		logarithm_table[365] = 14'b0000001_1000010;
		logarithm_table[366] = 14'b0000001_1000010;
		logarithm_table[367] = 14'b0000001_1000011;
		logarithm_table[368] = 14'b0000001_1000011;
		logarithm_table[369] = 14'b0000001_1000100;
		logarithm_table[370] = 14'b0000001_1000100;
		logarithm_table[371] = 14'b0000001_1000101;
		logarithm_table[372] = 14'b0000001_1000101;
		logarithm_table[373] = 14'b0000001_1000110;
		logarithm_table[374] = 14'b0000001_1000110;
		logarithm_table[375] = 14'b0000001_1000110;
		logarithm_table[376] = 14'b0000001_1000111;
		logarithm_table[377] = 14'b0000001_1000111;
		logarithm_table[378] = 14'b0000001_1001000;
		logarithm_table[379] = 14'b0000001_1001000;
		logarithm_table[380] = 14'b0000001_1001001;
		logarithm_table[381] = 14'b0000001_1001001;
		logarithm_table[382] = 14'b0000001_1001010;
		logarithm_table[383] = 14'b0000001_1001010;
		logarithm_table[384] = 14'b0000001_1001011;
		logarithm_table[385] = 14'b0000001_1001011;
		logarithm_table[386] = 14'b0000001_1001100;
		logarithm_table[387] = 14'b0000001_1001100;
		logarithm_table[388] = 14'b0000001_1001101;
		logarithm_table[389] = 14'b0000001_1001101;
		logarithm_table[390] = 14'b0000001_1001110;
		logarithm_table[391] = 14'b0000001_1001110;
		logarithm_table[392] = 14'b0000001_1001111;
		logarithm_table[393] = 14'b0000001_1001111;
		logarithm_table[394] = 14'b0000001_1010000;
		logarithm_table[395] = 14'b0000001_1010000;
		logarithm_table[396] = 14'b0000001_1010001;
		logarithm_table[397] = 14'b0000001_1010001;
		logarithm_table[398] = 14'b0000001_1010001;
		logarithm_table[399] = 14'b0000001_1010010;
		logarithm_table[400] = 14'b0000001_1010010;
		logarithm_table[401] = 14'b0000001_1010011;
		logarithm_table[402] = 14'b0000001_1010011;
		logarithm_table[403] = 14'b0000001_1010100;
		logarithm_table[404] = 14'b0000001_1010100;
		logarithm_table[405] = 14'b0000001_1010101;
		logarithm_table[406] = 14'b0000001_1010101;
		logarithm_table[407] = 14'b0000001_1010110;
		logarithm_table[408] = 14'b0000001_1010110;
		logarithm_table[409] = 14'b0000001_1010111;
		logarithm_table[410] = 14'b0000001_1010111;
		logarithm_table[411] = 14'b0000001_1010111;
		logarithm_table[412] = 14'b0000001_1011000;
		logarithm_table[413] = 14'b0000001_1011000;
		logarithm_table[414] = 14'b0000001_1011001;
		logarithm_table[415] = 14'b0000001_1011001;
		logarithm_table[416] = 14'b0000001_1011010;
		logarithm_table[417] = 14'b0000001_1011010;
		logarithm_table[418] = 14'b0000001_1011011;
		logarithm_table[419] = 14'b0000001_1011011;
		logarithm_table[420] = 14'b0000001_1011011;
		logarithm_table[421] = 14'b0000001_1011100;
		logarithm_table[422] = 14'b0000001_1011100;
		logarithm_table[423] = 14'b0000001_1011101;
		logarithm_table[424] = 14'b0000001_1011101;
		logarithm_table[425] = 14'b0000001_1011110;
		logarithm_table[426] = 14'b0000001_1011110;
		logarithm_table[427] = 14'b0000001_1011110;
		logarithm_table[428] = 14'b0000001_1011111;
		logarithm_table[429] = 14'b0000001_1011111;
		logarithm_table[430] = 14'b0000001_1100000;
		logarithm_table[431] = 14'b0000001_1100000;
		logarithm_table[432] = 14'b0000001_1100001;
		logarithm_table[433] = 14'b0000001_1100001;
		logarithm_table[434] = 14'b0000001_1100001;
		logarithm_table[435] = 14'b0000001_1100010;
		logarithm_table[436] = 14'b0000001_1100010;
		logarithm_table[437] = 14'b0000001_1100011;
		logarithm_table[438] = 14'b0000001_1100011;
		logarithm_table[439] = 14'b0000001_1100100;
		logarithm_table[440] = 14'b0000001_1100100;
		logarithm_table[441] = 14'b0000001_1100100;
		logarithm_table[442] = 14'b0000001_1100101;
		logarithm_table[443] = 14'b0000001_1100101;
		logarithm_table[444] = 14'b0000001_1100110;
		logarithm_table[445] = 14'b0000001_1100110;
		logarithm_table[446] = 14'b0000001_1100111;
		logarithm_table[447] = 14'b0000001_1100111;
		logarithm_table[448] = 14'b0000001_1100111;
		logarithm_table[449] = 14'b0000001_1101000;
		logarithm_table[450] = 14'b0000001_1101000;
		logarithm_table[451] = 14'b0000001_1101001;
		logarithm_table[452] = 14'b0000001_1101001;
		logarithm_table[453] = 14'b0000001_1101001;
		logarithm_table[454] = 14'b0000001_1101010;
		logarithm_table[455] = 14'b0000001_1101010;
		logarithm_table[456] = 14'b0000001_1101011;
		logarithm_table[457] = 14'b0000001_1101011;
		logarithm_table[458] = 14'b0000001_1101011;
		logarithm_table[459] = 14'b0000001_1101100;
		logarithm_table[460] = 14'b0000001_1101100;
		logarithm_table[461] = 14'b0000001_1101101;
		logarithm_table[462] = 14'b0000001_1101101;
		logarithm_table[463] = 14'b0000001_1101101;
		logarithm_table[464] = 14'b0000001_1101110;
		logarithm_table[465] = 14'b0000001_1101110;
		logarithm_table[466] = 14'b0000001_1101111;
		logarithm_table[467] = 14'b0000001_1101111;
		logarithm_table[468] = 14'b0000001_1101111;
		logarithm_table[469] = 14'b0000001_1110000;
		logarithm_table[470] = 14'b0000001_1110000;
		logarithm_table[471] = 14'b0000001_1110001;
		logarithm_table[472] = 14'b0000001_1110001;
		logarithm_table[473] = 14'b0000001_1110001;
		logarithm_table[474] = 14'b0000001_1110010;
		logarithm_table[475] = 14'b0000001_1110010;
		logarithm_table[476] = 14'b0000001_1110011;
		logarithm_table[477] = 14'b0000001_1110011;
		logarithm_table[478] = 14'b0000001_1110011;
		logarithm_table[479] = 14'b0000001_1110100;
		logarithm_table[480] = 14'b0000001_1110100;
		logarithm_table[481] = 14'b0000001_1110100;
		logarithm_table[482] = 14'b0000001_1110101;
		logarithm_table[483] = 14'b0000001_1110101;
		logarithm_table[484] = 14'b0000001_1110110;
		logarithm_table[485] = 14'b0000001_1110110;
		logarithm_table[486] = 14'b0000001_1110110;
		logarithm_table[487] = 14'b0000001_1110111;
		logarithm_table[488] = 14'b0000001_1110111;
		logarithm_table[489] = 14'b0000001_1111000;
		logarithm_table[490] = 14'b0000001_1111000;
		logarithm_table[491] = 14'b0000001_1111000;
		logarithm_table[492] = 14'b0000001_1111001;
		logarithm_table[493] = 14'b0000001_1111001;
		logarithm_table[494] = 14'b0000001_1111001;
		logarithm_table[495] = 14'b0000001_1111010;
		logarithm_table[496] = 14'b0000001_1111010;
		logarithm_table[497] = 14'b0000001_1111011;
		logarithm_table[498] = 14'b0000001_1111011;
		logarithm_table[499] = 14'b0000001_1111011;
		logarithm_table[500] = 14'b0000001_1111100;
		logarithm_table[501] = 14'b0000001_1111100;
		logarithm_table[502] = 14'b0000001_1111100;
		logarithm_table[503] = 14'b0000001_1111101;
		logarithm_table[504] = 14'b0000001_1111101;
		logarithm_table[505] = 14'b0000001_1111101;
		logarithm_table[506] = 14'b0000001_1111110;
		logarithm_table[507] = 14'b0000001_1111110;
		logarithm_table[508] = 14'b0000001_1111111;
		logarithm_table[509] = 14'b0000001_1111111;
		logarithm_table[510] = 14'b0000001_1111111;
		logarithm_table[511] = 14'b0000010_0000000;
		logarithm_table[512] = 14'b0000010_0000000;
		logarithm_table[513] = 14'b0000010_0000000;
		logarithm_table[514] = 14'b0000010_0000001;
		logarithm_table[515] = 14'b0000010_0000001;
		logarithm_table[516] = 14'b0000010_0000001;
		logarithm_table[517] = 14'b0000010_0000010;
		logarithm_table[518] = 14'b0000010_0000010;
		logarithm_table[519] = 14'b0000010_0000011;
		logarithm_table[520] = 14'b0000010_0000011;
		logarithm_table[521] = 14'b0000010_0000011;
		logarithm_table[522] = 14'b0000010_0000100;
		logarithm_table[523] = 14'b0000010_0000100;
		logarithm_table[524] = 14'b0000010_0000100;
		logarithm_table[525] = 14'b0000010_0000101;
		logarithm_table[526] = 14'b0000010_0000101;
		logarithm_table[527] = 14'b0000010_0000101;
		logarithm_table[528] = 14'b0000010_0000110;
		logarithm_table[529] = 14'b0000010_0000110;
		logarithm_table[530] = 14'b0000010_0000110;
		logarithm_table[531] = 14'b0000010_0000111;
		logarithm_table[532] = 14'b0000010_0000111;
		logarithm_table[533] = 14'b0000010_0000111;
		logarithm_table[534] = 14'b0000010_0001000;
		logarithm_table[535] = 14'b0000010_0001000;
		logarithm_table[536] = 14'b0000010_0001000;
		logarithm_table[537] = 14'b0000010_0001001;
		logarithm_table[538] = 14'b0000010_0001001;
		logarithm_table[539] = 14'b0000010_0001001;
		logarithm_table[540] = 14'b0000010_0001010;
		logarithm_table[541] = 14'b0000010_0001010;
		logarithm_table[542] = 14'b0000010_0001011;
		logarithm_table[543] = 14'b0000010_0001011;
		logarithm_table[544] = 14'b0000010_0001011;
		logarithm_table[545] = 14'b0000010_0001100;
		logarithm_table[546] = 14'b0000010_0001100;
		logarithm_table[547] = 14'b0000010_0001100;
		logarithm_table[548] = 14'b0000010_0001101;
		logarithm_table[549] = 14'b0000010_0001101;
		logarithm_table[550] = 14'b0000010_0001101;
		logarithm_table[551] = 14'b0000010_0001110;
		logarithm_table[552] = 14'b0000010_0001110;
		logarithm_table[553] = 14'b0000010_0001110;
		logarithm_table[554] = 14'b0000010_0001111;
		logarithm_table[555] = 14'b0000010_0001111;
		logarithm_table[556] = 14'b0000010_0001111;
		logarithm_table[557] = 14'b0000010_0010000;
		logarithm_table[558] = 14'b0000010_0010000;
		logarithm_table[559] = 14'b0000010_0010000;
		logarithm_table[560] = 14'b0000010_0010001;
		logarithm_table[561] = 14'b0000010_0010001;
		logarithm_table[562] = 14'b0000010_0010001;
		logarithm_table[563] = 14'b0000010_0010010;
		logarithm_table[564] = 14'b0000010_0010010;
		logarithm_table[565] = 14'b0000010_0010010;
		logarithm_table[566] = 14'b0000010_0010011;
		logarithm_table[567] = 14'b0000010_0010011;
		logarithm_table[568] = 14'b0000010_0010011;
		logarithm_table[569] = 14'b0000010_0010011;
		logarithm_table[570] = 14'b0000010_0010100;
		logarithm_table[571] = 14'b0000010_0010100;
		logarithm_table[572] = 14'b0000010_0010100;
		logarithm_table[573] = 14'b0000010_0010101;
		logarithm_table[574] = 14'b0000010_0010101;
		logarithm_table[575] = 14'b0000010_0010101;
		logarithm_table[576] = 14'b0000010_0010110;
		logarithm_table[577] = 14'b0000010_0010110;
		logarithm_table[578] = 14'b0000010_0010110;
		logarithm_table[579] = 14'b0000010_0010111;
		logarithm_table[580] = 14'b0000010_0010111;
		logarithm_table[581] = 14'b0000010_0010111;
		logarithm_table[582] = 14'b0000010_0011000;
		logarithm_table[583] = 14'b0000010_0011000;
		logarithm_table[584] = 14'b0000010_0011000;
		logarithm_table[585] = 14'b0000010_0011001;
		logarithm_table[586] = 14'b0000010_0011001;
		logarithm_table[587] = 14'b0000010_0011001;
		logarithm_table[588] = 14'b0000010_0011010;
		logarithm_table[589] = 14'b0000010_0011010;
		logarithm_table[590] = 14'b0000010_0011010;
		logarithm_table[591] = 14'b0000010_0011010;
		logarithm_table[592] = 14'b0000010_0011011;
		logarithm_table[593] = 14'b0000010_0011011;
		logarithm_table[594] = 14'b0000010_0011011;
		logarithm_table[595] = 14'b0000010_0011100;
		logarithm_table[596] = 14'b0000010_0011100;
		logarithm_table[597] = 14'b0000010_0011100;
		logarithm_table[598] = 14'b0000010_0011101;
		logarithm_table[599] = 14'b0000010_0011101;
		logarithm_table[600] = 14'b0000010_0011101;
		logarithm_table[601] = 14'b0000010_0011110;
		logarithm_table[602] = 14'b0000010_0011110;
		logarithm_table[603] = 14'b0000010_0011110;
		logarithm_table[604] = 14'b0000010_0011111;
		logarithm_table[605] = 14'b0000010_0011111;
		logarithm_table[606] = 14'b0000010_0011111;
		logarithm_table[607] = 14'b0000010_0011111;
		logarithm_table[608] = 14'b0000010_0100000;
		logarithm_table[609] = 14'b0000010_0100000;
		logarithm_table[610] = 14'b0000010_0100000;
		logarithm_table[611] = 14'b0000010_0100001;
		logarithm_table[612] = 14'b0000010_0100001;
		logarithm_table[613] = 14'b0000010_0100001;
		logarithm_table[614] = 14'b0000010_0100010;
		logarithm_table[615] = 14'b0000010_0100010;
		logarithm_table[616] = 14'b0000010_0100010;
		logarithm_table[617] = 14'b0000010_0100010;
		logarithm_table[618] = 14'b0000010_0100011;
		logarithm_table[619] = 14'b0000010_0100011;
		logarithm_table[620] = 14'b0000010_0100011;
		logarithm_table[621] = 14'b0000010_0100100;
		logarithm_table[622] = 14'b0000010_0100100;
		logarithm_table[623] = 14'b0000010_0100100;
		logarithm_table[624] = 14'b0000010_0100101;
		logarithm_table[625] = 14'b0000010_0100101;
		logarithm_table[626] = 14'b0000010_0100101;
		logarithm_table[627] = 14'b0000010_0100101;
		logarithm_table[628] = 14'b0000010_0100110;
		logarithm_table[629] = 14'b0000010_0100110;
		logarithm_table[630] = 14'b0000010_0100110;
		logarithm_table[631] = 14'b0000010_0100111;
		logarithm_table[632] = 14'b0000010_0100111;
		logarithm_table[633] = 14'b0000010_0100111;
		logarithm_table[634] = 14'b0000010_0100111;
		logarithm_table[635] = 14'b0000010_0101000;
		logarithm_table[636] = 14'b0000010_0101000;
		logarithm_table[637] = 14'b0000010_0101000;
		logarithm_table[638] = 14'b0000010_0101001;
		logarithm_table[639] = 14'b0000010_0101001;
		logarithm_table[640] = 14'b0000010_0101001;
		logarithm_table[641] = 14'b0000010_0101001;
		logarithm_table[642] = 14'b0000010_0101010;
		logarithm_table[643] = 14'b0000010_0101010;
		logarithm_table[644] = 14'b0000010_0101010;
		logarithm_table[645] = 14'b0000010_0101011;
		logarithm_table[646] = 14'b0000010_0101011;
		logarithm_table[647] = 14'b0000010_0101011;
		logarithm_table[648] = 14'b0000010_0101100;
		logarithm_table[649] = 14'b0000010_0101100;
		logarithm_table[650] = 14'b0000010_0101100;
		logarithm_table[651] = 14'b0000010_0101100;
		logarithm_table[652] = 14'b0000010_0101101;
		logarithm_table[653] = 14'b0000010_0101101;
		logarithm_table[654] = 14'b0000010_0101101;
		logarithm_table[655] = 14'b0000010_0101101;
		logarithm_table[656] = 14'b0000010_0101110;
		logarithm_table[657] = 14'b0000010_0101110;
		logarithm_table[658] = 14'b0000010_0101110;
		logarithm_table[659] = 14'b0000010_0101111;
		logarithm_table[660] = 14'b0000010_0101111;
		logarithm_table[661] = 14'b0000010_0101111;
		logarithm_table[662] = 14'b0000010_0101111;
		logarithm_table[663] = 14'b0000010_0110000;
		logarithm_table[664] = 14'b0000010_0110000;
		logarithm_table[665] = 14'b0000010_0110000;
		logarithm_table[666] = 14'b0000010_0110001;
		logarithm_table[667] = 14'b0000010_0110001;
		logarithm_table[668] = 14'b0000010_0110001;
		logarithm_table[669] = 14'b0000010_0110001;
		logarithm_table[670] = 14'b0000010_0110010;
		logarithm_table[671] = 14'b0000010_0110010;
		logarithm_table[672] = 14'b0000010_0110010;
		logarithm_table[673] = 14'b0000010_0110010;
		logarithm_table[674] = 14'b0000010_0110011;
		logarithm_table[675] = 14'b0000010_0110011;
		logarithm_table[676] = 14'b0000010_0110011;
		logarithm_table[677] = 14'b0000010_0110100;
		logarithm_table[678] = 14'b0000010_0110100;
		logarithm_table[679] = 14'b0000010_0110100;
		logarithm_table[680] = 14'b0000010_0110100;
		logarithm_table[681] = 14'b0000010_0110101;
		logarithm_table[682] = 14'b0000010_0110101;
		logarithm_table[683] = 14'b0000010_0110101;
		logarithm_table[684] = 14'b0000010_0110101;
		logarithm_table[685] = 14'b0000010_0110110;
		logarithm_table[686] = 14'b0000010_0110110;
		logarithm_table[687] = 14'b0000010_0110110;
		logarithm_table[688] = 14'b0000010_0110111;
		logarithm_table[689] = 14'b0000010_0110111;
		logarithm_table[690] = 14'b0000010_0110111;
		logarithm_table[691] = 14'b0000010_0110111;
		logarithm_table[692] = 14'b0000010_0111000;
		logarithm_table[693] = 14'b0000010_0111000;
		logarithm_table[694] = 14'b0000010_0111000;
		logarithm_table[695] = 14'b0000010_0111000;
		logarithm_table[696] = 14'b0000010_0111001;
		logarithm_table[697] = 14'b0000010_0111001;
		logarithm_table[698] = 14'b0000010_0111001;
		logarithm_table[699] = 14'b0000010_0111001;
		logarithm_table[700] = 14'b0000010_0111010;
		logarithm_table[701] = 14'b0000010_0111010;
		logarithm_table[702] = 14'b0000010_0111010;
		logarithm_table[703] = 14'b0000010_0111011;
		logarithm_table[704] = 14'b0000010_0111011;
		logarithm_table[705] = 14'b0000010_0111011;
		logarithm_table[706] = 14'b0000010_0111011;
		logarithm_table[707] = 14'b0000010_0111100;
		logarithm_table[708] = 14'b0000010_0111100;
		logarithm_table[709] = 14'b0000010_0111100;
		logarithm_table[710] = 14'b0000010_0111100;
		logarithm_table[711] = 14'b0000010_0111101;
		logarithm_table[712] = 14'b0000010_0111101;
		logarithm_table[713] = 14'b0000010_0111101;
		logarithm_table[714] = 14'b0000010_0111101;
		logarithm_table[715] = 14'b0000010_0111110;
		logarithm_table[716] = 14'b0000010_0111110;
		logarithm_table[717] = 14'b0000010_0111110;
		logarithm_table[718] = 14'b0000010_0111110;
		logarithm_table[719] = 14'b0000010_0111111;
		logarithm_table[720] = 14'b0000010_0111111;
		logarithm_table[721] = 14'b0000010_0111111;
		logarithm_table[722] = 14'b0000010_0111111;
		logarithm_table[723] = 14'b0000010_1000000;
		logarithm_table[724] = 14'b0000010_1000000;
		logarithm_table[725] = 14'b0000010_1000000;
		logarithm_table[726] = 14'b0000010_1000000;
		logarithm_table[727] = 14'b0000010_1000001;
		logarithm_table[728] = 14'b0000010_1000001;
		logarithm_table[729] = 14'b0000010_1000001;
		logarithm_table[730] = 14'b0000010_1000010;
		logarithm_table[731] = 14'b0000010_1000010;
		logarithm_table[732] = 14'b0000010_1000010;
		logarithm_table[733] = 14'b0000010_1000010;
		logarithm_table[734] = 14'b0000010_1000011;
		logarithm_table[735] = 14'b0000010_1000011;
		logarithm_table[736] = 14'b0000010_1000011;
		logarithm_table[737] = 14'b0000010_1000011;
		logarithm_table[738] = 14'b0000010_1000100;
		logarithm_table[739] = 14'b0000010_1000100;
		logarithm_table[740] = 14'b0000010_1000100;
		logarithm_table[741] = 14'b0000010_1000100;
		logarithm_table[742] = 14'b0000010_1000101;
		logarithm_table[743] = 14'b0000010_1000101;
		logarithm_table[744] = 14'b0000010_1000101;
		logarithm_table[745] = 14'b0000010_1000101;
		logarithm_table[746] = 14'b0000010_1000110;
		logarithm_table[747] = 14'b0000010_1000110;
		logarithm_table[748] = 14'b0000010_1000110;
		logarithm_table[749] = 14'b0000010_1000110;
		logarithm_table[750] = 14'b0000010_1000110;
		logarithm_table[751] = 14'b0000010_1000111;
		logarithm_table[752] = 14'b0000010_1000111;
		logarithm_table[753] = 14'b0000010_1000111;
		logarithm_table[754] = 14'b0000010_1000111;
		logarithm_table[755] = 14'b0000010_1001000;
		logarithm_table[756] = 14'b0000010_1001000;
		logarithm_table[757] = 14'b0000010_1001000;
		logarithm_table[758] = 14'b0000010_1001000;
		logarithm_table[759] = 14'b0000010_1001001;
		logarithm_table[760] = 14'b0000010_1001001;
		logarithm_table[761] = 14'b0000010_1001001;
		logarithm_table[762] = 14'b0000010_1001001;
		logarithm_table[763] = 14'b0000010_1001010;
		logarithm_table[764] = 14'b0000010_1001010;
		logarithm_table[765] = 14'b0000010_1001010;
		logarithm_table[766] = 14'b0000010_1001010;
		logarithm_table[767] = 14'b0000010_1001011;
		logarithm_table[768] = 14'b0000010_1001011;
		logarithm_table[769] = 14'b0000010_1001011;
		logarithm_table[770] = 14'b0000010_1001011;
		logarithm_table[771] = 14'b0000010_1001100;
		logarithm_table[772] = 14'b0000010_1001100;
		logarithm_table[773] = 14'b0000010_1001100;
		logarithm_table[774] = 14'b0000010_1001100;
		logarithm_table[775] = 14'b0000010_1001101;
		logarithm_table[776] = 14'b0000010_1001101;
		logarithm_table[777] = 14'b0000010_1001101;
		logarithm_table[778] = 14'b0000010_1001101;
		logarithm_table[779] = 14'b0000010_1001110;
		logarithm_table[780] = 14'b0000010_1001110;
		logarithm_table[781] = 14'b0000010_1001110;
		logarithm_table[782] = 14'b0000010_1001110;
		logarithm_table[783] = 14'b0000010_1001110;
		logarithm_table[784] = 14'b0000010_1001111;
		logarithm_table[785] = 14'b0000010_1001111;
		logarithm_table[786] = 14'b0000010_1001111;
		logarithm_table[787] = 14'b0000010_1001111;
		logarithm_table[788] = 14'b0000010_1010000;
		logarithm_table[789] = 14'b0000010_1010000;
		logarithm_table[790] = 14'b0000010_1010000;
		logarithm_table[791] = 14'b0000010_1010000;
		logarithm_table[792] = 14'b0000010_1010001;
		logarithm_table[793] = 14'b0000010_1010001;
		logarithm_table[794] = 14'b0000010_1010001;
		logarithm_table[795] = 14'b0000010_1010001;
		logarithm_table[796] = 14'b0000010_1010001;
		logarithm_table[797] = 14'b0000010_1010010;
		logarithm_table[798] = 14'b0000010_1010010;
		logarithm_table[799] = 14'b0000010_1010010;
		logarithm_table[800] = 14'b0000010_1010010;
		logarithm_table[801] = 14'b0000010_1010011;
		logarithm_table[802] = 14'b0000010_1010011;
		logarithm_table[803] = 14'b0000010_1010011;
		logarithm_table[804] = 14'b0000010_1010011;
		logarithm_table[805] = 14'b0000010_1010100;
		logarithm_table[806] = 14'b0000010_1010100;
		logarithm_table[807] = 14'b0000010_1010100;
		logarithm_table[808] = 14'b0000010_1010100;
		logarithm_table[809] = 14'b0000010_1010100;
		logarithm_table[810] = 14'b0000010_1010101;
		logarithm_table[811] = 14'b0000010_1010101;
		logarithm_table[812] = 14'b0000010_1010101;
		logarithm_table[813] = 14'b0000010_1010101;
		logarithm_table[814] = 14'b0000010_1010110;
		logarithm_table[815] = 14'b0000010_1010110;
		logarithm_table[816] = 14'b0000010_1010110;
		logarithm_table[817] = 14'b0000010_1010110;
		logarithm_table[818] = 14'b0000010_1010111;
		logarithm_table[819] = 14'b0000010_1010111;
		logarithm_table[820] = 14'b0000010_1010111;
		logarithm_table[821] = 14'b0000010_1010111;
		logarithm_table[822] = 14'b0000010_1010111;
		logarithm_table[823] = 14'b0000010_1011000;
		logarithm_table[824] = 14'b0000010_1011000;
		logarithm_table[825] = 14'b0000010_1011000;
		logarithm_table[826] = 14'b0000010_1011000;
		logarithm_table[827] = 14'b0000010_1011001;
		logarithm_table[828] = 14'b0000010_1011001;
		logarithm_table[829] = 14'b0000010_1011001;
		logarithm_table[830] = 14'b0000010_1011001;
		logarithm_table[831] = 14'b0000010_1011001;
		logarithm_table[832] = 14'b0000010_1011010;
		logarithm_table[833] = 14'b0000010_1011010;
		logarithm_table[834] = 14'b0000010_1011010;
		logarithm_table[835] = 14'b0000010_1011010;
		logarithm_table[836] = 14'b0000010_1011011;
		logarithm_table[837] = 14'b0000010_1011011;
		logarithm_table[838] = 14'b0000010_1011011;
		logarithm_table[839] = 14'b0000010_1011011;
		logarithm_table[840] = 14'b0000010_1011011;
		logarithm_table[841] = 14'b0000010_1011100;
		logarithm_table[842] = 14'b0000010_1011100;
		logarithm_table[843] = 14'b0000010_1011100;
		logarithm_table[844] = 14'b0000010_1011100;
		logarithm_table[845] = 14'b0000010_1011101;
		logarithm_table[846] = 14'b0000010_1011101;
		logarithm_table[847] = 14'b0000010_1011101;
		logarithm_table[848] = 14'b0000010_1011101;
		logarithm_table[849] = 14'b0000010_1011101;
		logarithm_table[850] = 14'b0000010_1011110;
		logarithm_table[851] = 14'b0000010_1011110;
		logarithm_table[852] = 14'b0000010_1011110;
		logarithm_table[853] = 14'b0000010_1011110;
		logarithm_table[854] = 14'b0000010_1011110;
		logarithm_table[855] = 14'b0000010_1011111;
		logarithm_table[856] = 14'b0000010_1011111;
		logarithm_table[857] = 14'b0000010_1011111;
		logarithm_table[858] = 14'b0000010_1011111;
		logarithm_table[859] = 14'b0000010_1100000;
		logarithm_table[860] = 14'b0000010_1100000;
		logarithm_table[861] = 14'b0000010_1100000;
		logarithm_table[862] = 14'b0000010_1100000;
		logarithm_table[863] = 14'b0000010_1100000;
		logarithm_table[864] = 14'b0000010_1100001;
		logarithm_table[865] = 14'b0000010_1100001;
		logarithm_table[866] = 14'b0000010_1100001;
		logarithm_table[867] = 14'b0000010_1100001;
		logarithm_table[868] = 14'b0000010_1100001;
		logarithm_table[869] = 14'b0000010_1100010;
		logarithm_table[870] = 14'b0000010_1100010;
		logarithm_table[871] = 14'b0000010_1100010;
		logarithm_table[872] = 14'b0000010_1100010;
		logarithm_table[873] = 14'b0000010_1100011;
		logarithm_table[874] = 14'b0000010_1100011;
		logarithm_table[875] = 14'b0000010_1100011;
		logarithm_table[876] = 14'b0000010_1100011;
		logarithm_table[877] = 14'b0000010_1100011;
		logarithm_table[878] = 14'b0000010_1100100;
		logarithm_table[879] = 14'b0000010_1100100;
		logarithm_table[880] = 14'b0000010_1100100;
		logarithm_table[881] = 14'b0000010_1100100;
		logarithm_table[882] = 14'b0000010_1100100;
		logarithm_table[883] = 14'b0000010_1100101;
		logarithm_table[884] = 14'b0000010_1100101;
		logarithm_table[885] = 14'b0000010_1100101;
		logarithm_table[886] = 14'b0000010_1100101;
		logarithm_table[887] = 14'b0000010_1100101;
		logarithm_table[888] = 14'b0000010_1100110;
		logarithm_table[889] = 14'b0000010_1100110;
		logarithm_table[890] = 14'b0000010_1100110;
		logarithm_table[891] = 14'b0000010_1100110;
		logarithm_table[892] = 14'b0000010_1100111;
		logarithm_table[893] = 14'b0000010_1100111;
		logarithm_table[894] = 14'b0000010_1100111;
		logarithm_table[895] = 14'b0000010_1100111;
		logarithm_table[896] = 14'b0000010_1100111;
		logarithm_table[897] = 14'b0000010_1101000;
		logarithm_table[898] = 14'b0000010_1101000;
		logarithm_table[899] = 14'b0000010_1101000;
		logarithm_table[900] = 14'b0000010_1101000;
		logarithm_table[901] = 14'b0000010_1101000;
		logarithm_table[902] = 14'b0000010_1101001;
		logarithm_table[903] = 14'b0000010_1101001;
		logarithm_table[904] = 14'b0000010_1101001;
		logarithm_table[905] = 14'b0000010_1101001;
		logarithm_table[906] = 14'b0000010_1101001;
		logarithm_table[907] = 14'b0000010_1101010;
		logarithm_table[908] = 14'b0000010_1101010;
		logarithm_table[909] = 14'b0000010_1101010;
		logarithm_table[910] = 14'b0000010_1101010;
		logarithm_table[911] = 14'b0000010_1101010;
		logarithm_table[912] = 14'b0000010_1101011;
		logarithm_table[913] = 14'b0000010_1101011;
		logarithm_table[914] = 14'b0000010_1101011;
		logarithm_table[915] = 14'b0000010_1101011;
		logarithm_table[916] = 14'b0000010_1101011;
		logarithm_table[917] = 14'b0000010_1101100;
		logarithm_table[918] = 14'b0000010_1101100;
		logarithm_table[919] = 14'b0000010_1101100;
		logarithm_table[920] = 14'b0000010_1101100;
		logarithm_table[921] = 14'b0000010_1101100;
		logarithm_table[922] = 14'b0000010_1101101;
		logarithm_table[923] = 14'b0000010_1101101;
		logarithm_table[924] = 14'b0000010_1101101;
		logarithm_table[925] = 14'b0000010_1101101;
		logarithm_table[926] = 14'b0000010_1101101;
		logarithm_table[927] = 14'b0000010_1101110;
		logarithm_table[928] = 14'b0000010_1101110;
		logarithm_table[929] = 14'b0000010_1101110;
		logarithm_table[930] = 14'b0000010_1101110;
		logarithm_table[931] = 14'b0000010_1101110;
		logarithm_table[932] = 14'b0000010_1101111;
		logarithm_table[933] = 14'b0000010_1101111;
		logarithm_table[934] = 14'b0000010_1101111;
		logarithm_table[935] = 14'b0000010_1101111;
		logarithm_table[936] = 14'b0000010_1101111;
		logarithm_table[937] = 14'b0000010_1110000;
		logarithm_table[938] = 14'b0000010_1110000;
		logarithm_table[939] = 14'b0000010_1110000;
		logarithm_table[940] = 14'b0000010_1110000;
		logarithm_table[941] = 14'b0000010_1110000;
		logarithm_table[942] = 14'b0000010_1110001;
		logarithm_table[943] = 14'b0000010_1110001;
		logarithm_table[944] = 14'b0000010_1110001;
		logarithm_table[945] = 14'b0000010_1110001;
		logarithm_table[946] = 14'b0000010_1110001;
		logarithm_table[947] = 14'b0000010_1110010;
		logarithm_table[948] = 14'b0000010_1110010;
		logarithm_table[949] = 14'b0000010_1110010;
		logarithm_table[950] = 14'b0000010_1110010;
		logarithm_table[951] = 14'b0000010_1110010;
		logarithm_table[952] = 14'b0000010_1110011;
		logarithm_table[953] = 14'b0000010_1110011;
		logarithm_table[954] = 14'b0000010_1110011;
		logarithm_table[955] = 14'b0000010_1110011;
		logarithm_table[956] = 14'b0000010_1110011;
		logarithm_table[957] = 14'b0000010_1110100;
		logarithm_table[958] = 14'b0000010_1110100;
		logarithm_table[959] = 14'b0000010_1110100;
		logarithm_table[960] = 14'b0000010_1110100;
		logarithm_table[961] = 14'b0000010_1110100;
		logarithm_table[962] = 14'b0000010_1110100;
		logarithm_table[963] = 14'b0000010_1110101;
		logarithm_table[964] = 14'b0000010_1110101;
		logarithm_table[965] = 14'b0000010_1110101;
		logarithm_table[966] = 14'b0000010_1110101;
		logarithm_table[967] = 14'b0000010_1110101;
		logarithm_table[968] = 14'b0000010_1110110;
		logarithm_table[969] = 14'b0000010_1110110;
		logarithm_table[970] = 14'b0000010_1110110;
		logarithm_table[971] = 14'b0000010_1110110;
		logarithm_table[972] = 14'b0000010_1110110;
		logarithm_table[973] = 14'b0000010_1110111;
		logarithm_table[974] = 14'b0000010_1110111;
		logarithm_table[975] = 14'b0000010_1110111;
		logarithm_table[976] = 14'b0000010_1110111;
		logarithm_table[977] = 14'b0000010_1110111;
		logarithm_table[978] = 14'b0000010_1111000;
		logarithm_table[979] = 14'b0000010_1111000;
		logarithm_table[980] = 14'b0000010_1111000;
		logarithm_table[981] = 14'b0000010_1111000;
		logarithm_table[982] = 14'b0000010_1111000;
		logarithm_table[983] = 14'b0000010_1111000;
		logarithm_table[984] = 14'b0000010_1111001;
		logarithm_table[985] = 14'b0000010_1111001;
		logarithm_table[986] = 14'b0000010_1111001;
		logarithm_table[987] = 14'b0000010_1111001;
		logarithm_table[988] = 14'b0000010_1111001;
		logarithm_table[989] = 14'b0000010_1111010;
		logarithm_table[990] = 14'b0000010_1111010;
		logarithm_table[991] = 14'b0000010_1111010;
		logarithm_table[992] = 14'b0000010_1111010;
		logarithm_table[993] = 14'b0000010_1111010;
		logarithm_table[994] = 14'b0000010_1111011;
		logarithm_table[995] = 14'b0000010_1111011;
		logarithm_table[996] = 14'b0000010_1111011;
		logarithm_table[997] = 14'b0000010_1111011;
		logarithm_table[998] = 14'b0000010_1111011;
		logarithm_table[999] = 14'b0000010_1111011;
		logarithm_table[1000] = 14'b0000010_1111100;
		logarithm_table[1001] = 14'b0000010_1111100;
		logarithm_table[1002] = 14'b0000010_1111100;
		logarithm_table[1003] = 14'b0000010_1111100;
		logarithm_table[1004] = 14'b0000010_1111100;
		logarithm_table[1005] = 14'b0000010_1111101;
		logarithm_table[1006] = 14'b0000010_1111101;
		logarithm_table[1007] = 14'b0000010_1111101;
		logarithm_table[1008] = 14'b0000010_1111101;
		logarithm_table[1009] = 14'b0000010_1111101;
		logarithm_table[1010] = 14'b0000010_1111101;
		logarithm_table[1011] = 14'b0000010_1111110;
		logarithm_table[1012] = 14'b0000010_1111110;
		logarithm_table[1013] = 14'b0000010_1111110;
		logarithm_table[1014] = 14'b0000010_1111110;
		logarithm_table[1015] = 14'b0000010_1111110;
		logarithm_table[1016] = 14'b0000010_1111111;
		logarithm_table[1017] = 14'b0000010_1111111;
		logarithm_table[1018] = 14'b0000010_1111111;
		logarithm_table[1019] = 14'b0000010_1111111;
		logarithm_table[1020] = 14'b0000010_1111111;
		logarithm_table[1021] = 14'b0000010_1111111;
		logarithm_table[1022] = 14'b0000011_0000000;
		logarithm_table[1023] = 14'b0000011_0000000;
		logarithm_table[1024] = 14'b0000011_0000000;
		logarithm_table[1025] = 14'b0000011_0000000;
		logarithm_table[1026] = 14'b0000011_0000000;
		logarithm_table[1027] = 14'b0000011_0000001;
		logarithm_table[1028] = 14'b0000011_0000001;
		logarithm_table[1029] = 14'b0000011_0000001;
		logarithm_table[1030] = 14'b0000011_0000001;
		logarithm_table[1031] = 14'b0000011_0000001;
		logarithm_table[1032] = 14'b0000011_0000001;
		logarithm_table[1033] = 14'b0000011_0000010;
		logarithm_table[1034] = 14'b0000011_0000010;
		logarithm_table[1035] = 14'b0000011_0000010;
		logarithm_table[1036] = 14'b0000011_0000010;
		logarithm_table[1037] = 14'b0000011_0000010;
		logarithm_table[1038] = 14'b0000011_0000011;
		logarithm_table[1039] = 14'b0000011_0000011;
		logarithm_table[1040] = 14'b0000011_0000011;
		logarithm_table[1041] = 14'b0000011_0000011;
		logarithm_table[1042] = 14'b0000011_0000011;
		logarithm_table[1043] = 14'b0000011_0000011;
		logarithm_table[1044] = 14'b0000011_0000100;
		logarithm_table[1045] = 14'b0000011_0000100;
		logarithm_table[1046] = 14'b0000011_0000100;
		logarithm_table[1047] = 14'b0000011_0000100;
		logarithm_table[1048] = 14'b0000011_0000100;
		logarithm_table[1049] = 14'b0000011_0000100;
		logarithm_table[1050] = 14'b0000011_0000101;
		logarithm_table[1051] = 14'b0000011_0000101;
		logarithm_table[1052] = 14'b0000011_0000101;
		logarithm_table[1053] = 14'b0000011_0000101;
		logarithm_table[1054] = 14'b0000011_0000101;
		logarithm_table[1055] = 14'b0000011_0000110;
		logarithm_table[1056] = 14'b0000011_0000110;
		logarithm_table[1057] = 14'b0000011_0000110;
		logarithm_table[1058] = 14'b0000011_0000110;
		logarithm_table[1059] = 14'b0000011_0000110;
		logarithm_table[1060] = 14'b0000011_0000110;
		logarithm_table[1061] = 14'b0000011_0000111;
		logarithm_table[1062] = 14'b0000011_0000111;
		logarithm_table[1063] = 14'b0000011_0000111;
		logarithm_table[1064] = 14'b0000011_0000111;
		logarithm_table[1065] = 14'b0000011_0000111;
		logarithm_table[1066] = 14'b0000011_0000111;
		logarithm_table[1067] = 14'b0000011_0001000;
		logarithm_table[1068] = 14'b0000011_0001000;
		logarithm_table[1069] = 14'b0000011_0001000;
		logarithm_table[1070] = 14'b0000011_0001000;
		logarithm_table[1071] = 14'b0000011_0001000;
		logarithm_table[1072] = 14'b0000011_0001000;
		logarithm_table[1073] = 14'b0000011_0001001;
		logarithm_table[1074] = 14'b0000011_0001001;
		logarithm_table[1075] = 14'b0000011_0001001;
		logarithm_table[1076] = 14'b0000011_0001001;
		logarithm_table[1077] = 14'b0000011_0001001;
		logarithm_table[1078] = 14'b0000011_0001001;
		logarithm_table[1079] = 14'b0000011_0001010;
		logarithm_table[1080] = 14'b0000011_0001010;
		logarithm_table[1081] = 14'b0000011_0001010;
		logarithm_table[1082] = 14'b0000011_0001010;
		logarithm_table[1083] = 14'b0000011_0001010;
		logarithm_table[1084] = 14'b0000011_0001011;
		logarithm_table[1085] = 14'b0000011_0001011;
		logarithm_table[1086] = 14'b0000011_0001011;
		logarithm_table[1087] = 14'b0000011_0001011;
		logarithm_table[1088] = 14'b0000011_0001011;
		logarithm_table[1089] = 14'b0000011_0001011;
		logarithm_table[1090] = 14'b0000011_0001100;
		logarithm_table[1091] = 14'b0000011_0001100;
		logarithm_table[1092] = 14'b0000011_0001100;
		logarithm_table[1093] = 14'b0000011_0001100;
		logarithm_table[1094] = 14'b0000011_0001100;
		logarithm_table[1095] = 14'b0000011_0001100;
		logarithm_table[1096] = 14'b0000011_0001101;
		logarithm_table[1097] = 14'b0000011_0001101;
		logarithm_table[1098] = 14'b0000011_0001101;
		logarithm_table[1099] = 14'b0000011_0001101;
		logarithm_table[1100] = 14'b0000011_0001101;
		logarithm_table[1101] = 14'b0000011_0001101;
		logarithm_table[1102] = 14'b0000011_0001110;
		logarithm_table[1103] = 14'b0000011_0001110;
		logarithm_table[1104] = 14'b0000011_0001110;
		logarithm_table[1105] = 14'b0000011_0001110;
		logarithm_table[1106] = 14'b0000011_0001110;
		logarithm_table[1107] = 14'b0000011_0001110;
		logarithm_table[1108] = 14'b0000011_0001111;
		logarithm_table[1109] = 14'b0000011_0001111;
		logarithm_table[1110] = 14'b0000011_0001111;
		logarithm_table[1111] = 14'b0000011_0001111;
		logarithm_table[1112] = 14'b0000011_0001111;
		logarithm_table[1113] = 14'b0000011_0001111;
		logarithm_table[1114] = 14'b0000011_0010000;
		logarithm_table[1115] = 14'b0000011_0010000;
		logarithm_table[1116] = 14'b0000011_0010000;
		logarithm_table[1117] = 14'b0000011_0010000;
		logarithm_table[1118] = 14'b0000011_0010000;
		logarithm_table[1119] = 14'b0000011_0010000;
		logarithm_table[1120] = 14'b0000011_0010001;
		logarithm_table[1121] = 14'b0000011_0010001;
		logarithm_table[1122] = 14'b0000011_0010001;
		logarithm_table[1123] = 14'b0000011_0010001;
		logarithm_table[1124] = 14'b0000011_0010001;
		logarithm_table[1125] = 14'b0000011_0010001;
		logarithm_table[1126] = 14'b0000011_0010010;
		logarithm_table[1127] = 14'b0000011_0010010;
		logarithm_table[1128] = 14'b0000011_0010010;
		logarithm_table[1129] = 14'b0000011_0010010;
		logarithm_table[1130] = 14'b0000011_0010010;
		logarithm_table[1131] = 14'b0000011_0010010;
		logarithm_table[1132] = 14'b0000011_0010011;
		logarithm_table[1133] = 14'b0000011_0010011;
		logarithm_table[1134] = 14'b0000011_0010011;
		logarithm_table[1135] = 14'b0000011_0010011;
		logarithm_table[1136] = 14'b0000011_0010011;
		logarithm_table[1137] = 14'b0000011_0010011;
		logarithm_table[1138] = 14'b0000011_0010011;
		logarithm_table[1139] = 14'b0000011_0010100;
		logarithm_table[1140] = 14'b0000011_0010100;
		logarithm_table[1141] = 14'b0000011_0010100;
		logarithm_table[1142] = 14'b0000011_0010100;
		logarithm_table[1143] = 14'b0000011_0010100;
		logarithm_table[1144] = 14'b0000011_0010100;
		logarithm_table[1145] = 14'b0000011_0010101;
		logarithm_table[1146] = 14'b0000011_0010101;
		logarithm_table[1147] = 14'b0000011_0010101;
		logarithm_table[1148] = 14'b0000011_0010101;
		logarithm_table[1149] = 14'b0000011_0010101;
		logarithm_table[1150] = 14'b0000011_0010101;
		logarithm_table[1151] = 14'b0000011_0010110;
		logarithm_table[1152] = 14'b0000011_0010110;
		logarithm_table[1153] = 14'b0000011_0010110;
		logarithm_table[1154] = 14'b0000011_0010110;
		logarithm_table[1155] = 14'b0000011_0010110;
		logarithm_table[1156] = 14'b0000011_0010110;
		logarithm_table[1157] = 14'b0000011_0010111;
		logarithm_table[1158] = 14'b0000011_0010111;
		logarithm_table[1159] = 14'b0000011_0010111;
		logarithm_table[1160] = 14'b0000011_0010111;
		logarithm_table[1161] = 14'b0000011_0010111;
		logarithm_table[1162] = 14'b0000011_0010111;
		logarithm_table[1163] = 14'b0000011_0011000;
		logarithm_table[1164] = 14'b0000011_0011000;
		logarithm_table[1165] = 14'b0000011_0011000;
		logarithm_table[1166] = 14'b0000011_0011000;
		logarithm_table[1167] = 14'b0000011_0011000;
		logarithm_table[1168] = 14'b0000011_0011000;
		logarithm_table[1169] = 14'b0000011_0011000;
		logarithm_table[1170] = 14'b0000011_0011001;
		logarithm_table[1171] = 14'b0000011_0011001;
		logarithm_table[1172] = 14'b0000011_0011001;
		logarithm_table[1173] = 14'b0000011_0011001;
		logarithm_table[1174] = 14'b0000011_0011001;
		logarithm_table[1175] = 14'b0000011_0011001;
		logarithm_table[1176] = 14'b0000011_0011010;
		logarithm_table[1177] = 14'b0000011_0011010;
		logarithm_table[1178] = 14'b0000011_0011010;
		logarithm_table[1179] = 14'b0000011_0011010;
		logarithm_table[1180] = 14'b0000011_0011010;
		logarithm_table[1181] = 14'b0000011_0011010;
		logarithm_table[1182] = 14'b0000011_0011010;
		logarithm_table[1183] = 14'b0000011_0011011;
		logarithm_table[1184] = 14'b0000011_0011011;
		logarithm_table[1185] = 14'b0000011_0011011;
		logarithm_table[1186] = 14'b0000011_0011011;
		logarithm_table[1187] = 14'b0000011_0011011;
		logarithm_table[1188] = 14'b0000011_0011011;
		logarithm_table[1189] = 14'b0000011_0011100;
		logarithm_table[1190] = 14'b0000011_0011100;
		logarithm_table[1191] = 14'b0000011_0011100;
		logarithm_table[1192] = 14'b0000011_0011100;
		logarithm_table[1193] = 14'b0000011_0011100;
		logarithm_table[1194] = 14'b0000011_0011100;
		logarithm_table[1195] = 14'b0000011_0011101;
		logarithm_table[1196] = 14'b0000011_0011101;
		logarithm_table[1197] = 14'b0000011_0011101;
		logarithm_table[1198] = 14'b0000011_0011101;
		logarithm_table[1199] = 14'b0000011_0011101;
		logarithm_table[1200] = 14'b0000011_0011101;
		logarithm_table[1201] = 14'b0000011_0011101;
		logarithm_table[1202] = 14'b0000011_0011110;
		logarithm_table[1203] = 14'b0000011_0011110;
		logarithm_table[1204] = 14'b0000011_0011110;
		logarithm_table[1205] = 14'b0000011_0011110;
		logarithm_table[1206] = 14'b0000011_0011110;
		logarithm_table[1207] = 14'b0000011_0011110;
		logarithm_table[1208] = 14'b0000011_0011111;
		logarithm_table[1209] = 14'b0000011_0011111;
		logarithm_table[1210] = 14'b0000011_0011111;
		logarithm_table[1211] = 14'b0000011_0011111;
		logarithm_table[1212] = 14'b0000011_0011111;
		logarithm_table[1213] = 14'b0000011_0011111;
		logarithm_table[1214] = 14'b0000011_0011111;
		logarithm_table[1215] = 14'b0000011_0100000;
		logarithm_table[1216] = 14'b0000011_0100000;
		logarithm_table[1217] = 14'b0000011_0100000;
		logarithm_table[1218] = 14'b0000011_0100000;
		logarithm_table[1219] = 14'b0000011_0100000;
		logarithm_table[1220] = 14'b0000011_0100000;
		logarithm_table[1221] = 14'b0000011_0100000;
		logarithm_table[1222] = 14'b0000011_0100001;
		logarithm_table[1223] = 14'b0000011_0100001;
		logarithm_table[1224] = 14'b0000011_0100001;
		logarithm_table[1225] = 14'b0000011_0100001;
		logarithm_table[1226] = 14'b0000011_0100001;
		logarithm_table[1227] = 14'b0000011_0100001;
		logarithm_table[1228] = 14'b0000011_0100010;
		logarithm_table[1229] = 14'b0000011_0100010;
		logarithm_table[1230] = 14'b0000011_0100010;
		logarithm_table[1231] = 14'b0000011_0100010;
		logarithm_table[1232] = 14'b0000011_0100010;
		logarithm_table[1233] = 14'b0000011_0100010;
		logarithm_table[1234] = 14'b0000011_0100010;
		logarithm_table[1235] = 14'b0000011_0100011;
		logarithm_table[1236] = 14'b0000011_0100011;
		logarithm_table[1237] = 14'b0000011_0100011;
		logarithm_table[1238] = 14'b0000011_0100011;
		logarithm_table[1239] = 14'b0000011_0100011;
		logarithm_table[1240] = 14'b0000011_0100011;
		logarithm_table[1241] = 14'b0000011_0100011;
		logarithm_table[1242] = 14'b0000011_0100100;
		logarithm_table[1243] = 14'b0000011_0100100;
		logarithm_table[1244] = 14'b0000011_0100100;
		logarithm_table[1245] = 14'b0000011_0100100;
		logarithm_table[1246] = 14'b0000011_0100100;
		logarithm_table[1247] = 14'b0000011_0100100;
		logarithm_table[1248] = 14'b0000011_0100101;
		logarithm_table[1249] = 14'b0000011_0100101;
		logarithm_table[1250] = 14'b0000011_0100101;
		logarithm_table[1251] = 14'b0000011_0100101;
		logarithm_table[1252] = 14'b0000011_0100101;
		logarithm_table[1253] = 14'b0000011_0100101;
		logarithm_table[1254] = 14'b0000011_0100101;
		logarithm_table[1255] = 14'b0000011_0100110;
		logarithm_table[1256] = 14'b0000011_0100110;
		logarithm_table[1257] = 14'b0000011_0100110;
		logarithm_table[1258] = 14'b0000011_0100110;
		logarithm_table[1259] = 14'b0000011_0100110;
		logarithm_table[1260] = 14'b0000011_0100110;
		logarithm_table[1261] = 14'b0000011_0100110;
		logarithm_table[1262] = 14'b0000011_0100111;
		logarithm_table[1263] = 14'b0000011_0100111;
		logarithm_table[1264] = 14'b0000011_0100111;
		logarithm_table[1265] = 14'b0000011_0100111;
		logarithm_table[1266] = 14'b0000011_0100111;
		logarithm_table[1267] = 14'b0000011_0100111;
		logarithm_table[1268] = 14'b0000011_0100111;
		logarithm_table[1269] = 14'b0000011_0101000;
		logarithm_table[1270] = 14'b0000011_0101000;
		logarithm_table[1271] = 14'b0000011_0101000;
		logarithm_table[1272] = 14'b0000011_0101000;
		logarithm_table[1273] = 14'b0000011_0101000;
		logarithm_table[1274] = 14'b0000011_0101000;
		logarithm_table[1275] = 14'b0000011_0101000;
		logarithm_table[1276] = 14'b0000011_0101001;
		logarithm_table[1277] = 14'b0000011_0101001;
		logarithm_table[1278] = 14'b0000011_0101001;
		logarithm_table[1279] = 14'b0000011_0101001;
		logarithm_table[1280] = 14'b0000011_0101001;
		logarithm_table[1281] = 14'b0000011_0101001;
		logarithm_table[1282] = 14'b0000011_0101001;
		logarithm_table[1283] = 14'b0000011_0101010;
		logarithm_table[1284] = 14'b0000011_0101010;
		logarithm_table[1285] = 14'b0000011_0101010;
		logarithm_table[1286] = 14'b0000011_0101010;
		logarithm_table[1287] = 14'b0000011_0101010;
		logarithm_table[1288] = 14'b0000011_0101010;
		logarithm_table[1289] = 14'b0000011_0101011;
		logarithm_table[1290] = 14'b0000011_0101011;
		logarithm_table[1291] = 14'b0000011_0101011;
		logarithm_table[1292] = 14'b0000011_0101011;
		logarithm_table[1293] = 14'b0000011_0101011;
		logarithm_table[1294] = 14'b0000011_0101011;
		logarithm_table[1295] = 14'b0000011_0101011;
		logarithm_table[1296] = 14'b0000011_0101100;
		logarithm_table[1297] = 14'b0000011_0101100;
		logarithm_table[1298] = 14'b0000011_0101100;
		logarithm_table[1299] = 14'b0000011_0101100;
		logarithm_table[1300] = 14'b0000011_0101100;
		logarithm_table[1301] = 14'b0000011_0101100;
		logarithm_table[1302] = 14'b0000011_0101100;
		logarithm_table[1303] = 14'b0000011_0101100;
		logarithm_table[1304] = 14'b0000011_0101101;
		logarithm_table[1305] = 14'b0000011_0101101;
		logarithm_table[1306] = 14'b0000011_0101101;
		logarithm_table[1307] = 14'b0000011_0101101;
		logarithm_table[1308] = 14'b0000011_0101101;
		logarithm_table[1309] = 14'b0000011_0101101;
		logarithm_table[1310] = 14'b0000011_0101101;
		logarithm_table[1311] = 14'b0000011_0101110;
		logarithm_table[1312] = 14'b0000011_0101110;
		logarithm_table[1313] = 14'b0000011_0101110;
		logarithm_table[1314] = 14'b0000011_0101110;
		logarithm_table[1315] = 14'b0000011_0101110;
		logarithm_table[1316] = 14'b0000011_0101110;
		logarithm_table[1317] = 14'b0000011_0101110;
		logarithm_table[1318] = 14'b0000011_0101111;
		logarithm_table[1319] = 14'b0000011_0101111;
		logarithm_table[1320] = 14'b0000011_0101111;
		logarithm_table[1321] = 14'b0000011_0101111;
		logarithm_table[1322] = 14'b0000011_0101111;
		logarithm_table[1323] = 14'b0000011_0101111;
		logarithm_table[1324] = 14'b0000011_0101111;
		logarithm_table[1325] = 14'b0000011_0110000;
		logarithm_table[1326] = 14'b0000011_0110000;
		logarithm_table[1327] = 14'b0000011_0110000;
		logarithm_table[1328] = 14'b0000011_0110000;
		logarithm_table[1329] = 14'b0000011_0110000;
		logarithm_table[1330] = 14'b0000011_0110000;
		logarithm_table[1331] = 14'b0000011_0110000;
		logarithm_table[1332] = 14'b0000011_0110001;
		logarithm_table[1333] = 14'b0000011_0110001;
		logarithm_table[1334] = 14'b0000011_0110001;
		logarithm_table[1335] = 14'b0000011_0110001;
		logarithm_table[1336] = 14'b0000011_0110001;
		logarithm_table[1337] = 14'b0000011_0110001;
		logarithm_table[1338] = 14'b0000011_0110001;
		logarithm_table[1339] = 14'b0000011_0110010;
		logarithm_table[1340] = 14'b0000011_0110010;
		logarithm_table[1341] = 14'b0000011_0110010;
		logarithm_table[1342] = 14'b0000011_0110010;
		logarithm_table[1343] = 14'b0000011_0110010;
		logarithm_table[1344] = 14'b0000011_0110010;
		logarithm_table[1345] = 14'b0000011_0110010;
		logarithm_table[1346] = 14'b0000011_0110010;
		logarithm_table[1347] = 14'b0000011_0110011;
		logarithm_table[1348] = 14'b0000011_0110011;
		logarithm_table[1349] = 14'b0000011_0110011;
		logarithm_table[1350] = 14'b0000011_0110011;
		logarithm_table[1351] = 14'b0000011_0110011;
		logarithm_table[1352] = 14'b0000011_0110011;
		logarithm_table[1353] = 14'b0000011_0110011;
		logarithm_table[1354] = 14'b0000011_0110100;
		logarithm_table[1355] = 14'b0000011_0110100;
		logarithm_table[1356] = 14'b0000011_0110100;
		logarithm_table[1357] = 14'b0000011_0110100;
		logarithm_table[1358] = 14'b0000011_0110100;
		logarithm_table[1359] = 14'b0000011_0110100;
		logarithm_table[1360] = 14'b0000011_0110100;
		logarithm_table[1361] = 14'b0000011_0110101;
		logarithm_table[1362] = 14'b0000011_0110101;
		logarithm_table[1363] = 14'b0000011_0110101;
		logarithm_table[1364] = 14'b0000011_0110101;
		logarithm_table[1365] = 14'b0000011_0110101;
		logarithm_table[1366] = 14'b0000011_0110101;
		logarithm_table[1367] = 14'b0000011_0110101;
		logarithm_table[1368] = 14'b0000011_0110101;
		logarithm_table[1369] = 14'b0000011_0110110;
		logarithm_table[1370] = 14'b0000011_0110110;
		logarithm_table[1371] = 14'b0000011_0110110;
		logarithm_table[1372] = 14'b0000011_0110110;
		logarithm_table[1373] = 14'b0000011_0110110;
		logarithm_table[1374] = 14'b0000011_0110110;
		logarithm_table[1375] = 14'b0000011_0110110;
		logarithm_table[1376] = 14'b0000011_0110111;
		logarithm_table[1377] = 14'b0000011_0110111;
		logarithm_table[1378] = 14'b0000011_0110111;
		logarithm_table[1379] = 14'b0000011_0110111;
		logarithm_table[1380] = 14'b0000011_0110111;
		logarithm_table[1381] = 14'b0000011_0110111;
		logarithm_table[1382] = 14'b0000011_0110111;
		logarithm_table[1383] = 14'b0000011_0110111;
		logarithm_table[1384] = 14'b0000011_0111000;
		logarithm_table[1385] = 14'b0000011_0111000;
		logarithm_table[1386] = 14'b0000011_0111000;
		logarithm_table[1387] = 14'b0000011_0111000;
		logarithm_table[1388] = 14'b0000011_0111000;
		logarithm_table[1389] = 14'b0000011_0111000;
		logarithm_table[1390] = 14'b0000011_0111000;
		logarithm_table[1391] = 14'b0000011_0111001;
		logarithm_table[1392] = 14'b0000011_0111001;
		logarithm_table[1393] = 14'b0000011_0111001;
		logarithm_table[1394] = 14'b0000011_0111001;
		logarithm_table[1395] = 14'b0000011_0111001;
		logarithm_table[1396] = 14'b0000011_0111001;
		logarithm_table[1397] = 14'b0000011_0111001;
		logarithm_table[1398] = 14'b0000011_0111001;
		logarithm_table[1399] = 14'b0000011_0111010;
		logarithm_table[1400] = 14'b0000011_0111010;
		logarithm_table[1401] = 14'b0000011_0111010;
		logarithm_table[1402] = 14'b0000011_0111010;
		logarithm_table[1403] = 14'b0000011_0111010;
		logarithm_table[1404] = 14'b0000011_0111010;
		logarithm_table[1405] = 14'b0000011_0111010;
		logarithm_table[1406] = 14'b0000011_0111011;
		logarithm_table[1407] = 14'b0000011_0111011;
		logarithm_table[1408] = 14'b0000011_0111011;
		logarithm_table[1409] = 14'b0000011_0111011;
		logarithm_table[1410] = 14'b0000011_0111011;
		logarithm_table[1411] = 14'b0000011_0111011;
		logarithm_table[1412] = 14'b0000011_0111011;
		logarithm_table[1413] = 14'b0000011_0111011;
		logarithm_table[1414] = 14'b0000011_0111100;
		logarithm_table[1415] = 14'b0000011_0111100;
		logarithm_table[1416] = 14'b0000011_0111100;
		logarithm_table[1417] = 14'b0000011_0111100;
		logarithm_table[1418] = 14'b0000011_0111100;
		logarithm_table[1419] = 14'b0000011_0111100;
		logarithm_table[1420] = 14'b0000011_0111100;
		logarithm_table[1421] = 14'b0000011_0111101;
		logarithm_table[1422] = 14'b0000011_0111101;
		logarithm_table[1423] = 14'b0000011_0111101;
		logarithm_table[1424] = 14'b0000011_0111101;
		logarithm_table[1425] = 14'b0000011_0111101;
		logarithm_table[1426] = 14'b0000011_0111101;
		logarithm_table[1427] = 14'b0000011_0111101;
		logarithm_table[1428] = 14'b0000011_0111101;
		logarithm_table[1429] = 14'b0000011_0111110;
		logarithm_table[1430] = 14'b0000011_0111110;
		logarithm_table[1431] = 14'b0000011_0111110;
		logarithm_table[1432] = 14'b0000011_0111110;
		logarithm_table[1433] = 14'b0000011_0111110;
		logarithm_table[1434] = 14'b0000011_0111110;
		logarithm_table[1435] = 14'b0000011_0111110;
		logarithm_table[1436] = 14'b0000011_0111110;
		logarithm_table[1437] = 14'b0000011_0111111;
		logarithm_table[1438] = 14'b0000011_0111111;
		logarithm_table[1439] = 14'b0000011_0111111;
		logarithm_table[1440] = 14'b0000011_0111111;
		logarithm_table[1441] = 14'b0000011_0111111;
		logarithm_table[1442] = 14'b0000011_0111111;
		logarithm_table[1443] = 14'b0000011_0111111;
		logarithm_table[1444] = 14'b0000011_0111111;
		logarithm_table[1445] = 14'b0000011_1000000;
		logarithm_table[1446] = 14'b0000011_1000000;
		logarithm_table[1447] = 14'b0000011_1000000;
		logarithm_table[1448] = 14'b0000011_1000000;
		logarithm_table[1449] = 14'b0000011_1000000;
		logarithm_table[1450] = 14'b0000011_1000000;
		logarithm_table[1451] = 14'b0000011_1000000;
		logarithm_table[1452] = 14'b0000011_1000000;
		logarithm_table[1453] = 14'b0000011_1000001;
		logarithm_table[1454] = 14'b0000011_1000001;
		logarithm_table[1455] = 14'b0000011_1000001;
		logarithm_table[1456] = 14'b0000011_1000001;
		logarithm_table[1457] = 14'b0000011_1000001;
		logarithm_table[1458] = 14'b0000011_1000001;
		logarithm_table[1459] = 14'b0000011_1000001;
		logarithm_table[1460] = 14'b0000011_1000010;
		logarithm_table[1461] = 14'b0000011_1000010;
		logarithm_table[1462] = 14'b0000011_1000010;
		logarithm_table[1463] = 14'b0000011_1000010;
		logarithm_table[1464] = 14'b0000011_1000010;
		logarithm_table[1465] = 14'b0000011_1000010;
		logarithm_table[1466] = 14'b0000011_1000010;
		logarithm_table[1467] = 14'b0000011_1000010;
		logarithm_table[1468] = 14'b0000011_1000011;
		logarithm_table[1469] = 14'b0000011_1000011;
		logarithm_table[1470] = 14'b0000011_1000011;
		logarithm_table[1471] = 14'b0000011_1000011;
		logarithm_table[1472] = 14'b0000011_1000011;
		logarithm_table[1473] = 14'b0000011_1000011;
		logarithm_table[1474] = 14'b0000011_1000011;
		logarithm_table[1475] = 14'b0000011_1000011;
		logarithm_table[1476] = 14'b0000011_1000100;
		logarithm_table[1477] = 14'b0000011_1000100;
		logarithm_table[1478] = 14'b0000011_1000100;
		logarithm_table[1479] = 14'b0000011_1000100;
		logarithm_table[1480] = 14'b0000011_1000100;
		logarithm_table[1481] = 14'b0000011_1000100;
		logarithm_table[1482] = 14'b0000011_1000100;
		logarithm_table[1483] = 14'b0000011_1000100;
		logarithm_table[1484] = 14'b0000011_1000101;
		logarithm_table[1485] = 14'b0000011_1000101;
		logarithm_table[1486] = 14'b0000011_1000101;
		logarithm_table[1487] = 14'b0000011_1000101;
		logarithm_table[1488] = 14'b0000011_1000101;
		logarithm_table[1489] = 14'b0000011_1000101;
		logarithm_table[1490] = 14'b0000011_1000101;
		logarithm_table[1491] = 14'b0000011_1000101;
		logarithm_table[1492] = 14'b0000011_1000110;
		logarithm_table[1493] = 14'b0000011_1000110;
		logarithm_table[1494] = 14'b0000011_1000110;
		logarithm_table[1495] = 14'b0000011_1000110;
		logarithm_table[1496] = 14'b0000011_1000110;
		logarithm_table[1497] = 14'b0000011_1000110;
		logarithm_table[1498] = 14'b0000011_1000110;
		logarithm_table[1499] = 14'b0000011_1000110;
		logarithm_table[1500] = 14'b0000011_1000110;
		logarithm_table[1501] = 14'b0000011_1000111;
		logarithm_table[1502] = 14'b0000011_1000111;
		logarithm_table[1503] = 14'b0000011_1000111;
		logarithm_table[1504] = 14'b0000011_1000111;
		logarithm_table[1505] = 14'b0000011_1000111;
		logarithm_table[1506] = 14'b0000011_1000111;
		logarithm_table[1507] = 14'b0000011_1000111;
		logarithm_table[1508] = 14'b0000011_1000111;
		logarithm_table[1509] = 14'b0000011_1001000;
		logarithm_table[1510] = 14'b0000011_1001000;
		logarithm_table[1511] = 14'b0000011_1001000;
		logarithm_table[1512] = 14'b0000011_1001000;
		logarithm_table[1513] = 14'b0000011_1001000;
		logarithm_table[1514] = 14'b0000011_1001000;
		logarithm_table[1515] = 14'b0000011_1001000;
		logarithm_table[1516] = 14'b0000011_1001000;
		logarithm_table[1517] = 14'b0000011_1001001;
		logarithm_table[1518] = 14'b0000011_1001001;
		logarithm_table[1519] = 14'b0000011_1001001;
		logarithm_table[1520] = 14'b0000011_1001001;
		logarithm_table[1521] = 14'b0000011_1001001;
		logarithm_table[1522] = 14'b0000011_1001001;
		logarithm_table[1523] = 14'b0000011_1001001;
		logarithm_table[1524] = 14'b0000011_1001001;
		logarithm_table[1525] = 14'b0000011_1001010;
		logarithm_table[1526] = 14'b0000011_1001010;
		logarithm_table[1527] = 14'b0000011_1001010;
		logarithm_table[1528] = 14'b0000011_1001010;
		logarithm_table[1529] = 14'b0000011_1001010;
		logarithm_table[1530] = 14'b0000011_1001010;
		logarithm_table[1531] = 14'b0000011_1001010;
		logarithm_table[1532] = 14'b0000011_1001010;
		logarithm_table[1533] = 14'b0000011_1001011;
		logarithm_table[1534] = 14'b0000011_1001011;
		logarithm_table[1535] = 14'b0000011_1001011;
		logarithm_table[1536] = 14'b0000011_1001011;
		logarithm_table[1537] = 14'b0000011_1001011;
		logarithm_table[1538] = 14'b0000011_1001011;
		logarithm_table[1539] = 14'b0000011_1001011;
		logarithm_table[1540] = 14'b0000011_1001011;
		logarithm_table[1541] = 14'b0000011_1001011;
		logarithm_table[1542] = 14'b0000011_1001100;
		logarithm_table[1543] = 14'b0000011_1001100;
		logarithm_table[1544] = 14'b0000011_1001100;
		logarithm_table[1545] = 14'b0000011_1001100;
		logarithm_table[1546] = 14'b0000011_1001100;
		logarithm_table[1547] = 14'b0000011_1001100;
		logarithm_table[1548] = 14'b0000011_1001100;
		logarithm_table[1549] = 14'b0000011_1001100;
		logarithm_table[1550] = 14'b0000011_1001101;
		logarithm_table[1551] = 14'b0000011_1001101;
		logarithm_table[1552] = 14'b0000011_1001101;
		logarithm_table[1553] = 14'b0000011_1001101;
		logarithm_table[1554] = 14'b0000011_1001101;
		logarithm_table[1555] = 14'b0000011_1001101;
		logarithm_table[1556] = 14'b0000011_1001101;
		logarithm_table[1557] = 14'b0000011_1001101;
		logarithm_table[1558] = 14'b0000011_1001110;
		logarithm_table[1559] = 14'b0000011_1001110;
		logarithm_table[1560] = 14'b0000011_1001110;
		logarithm_table[1561] = 14'b0000011_1001110;
		logarithm_table[1562] = 14'b0000011_1001110;
		logarithm_table[1563] = 14'b0000011_1001110;
		logarithm_table[1564] = 14'b0000011_1001110;
		logarithm_table[1565] = 14'b0000011_1001110;
		logarithm_table[1566] = 14'b0000011_1001110;
		logarithm_table[1567] = 14'b0000011_1001111;
		logarithm_table[1568] = 14'b0000011_1001111;
		logarithm_table[1569] = 14'b0000011_1001111;
		logarithm_table[1570] = 14'b0000011_1001111;
		logarithm_table[1571] = 14'b0000011_1001111;
		logarithm_table[1572] = 14'b0000011_1001111;
		logarithm_table[1573] = 14'b0000011_1001111;
		logarithm_table[1574] = 14'b0000011_1001111;
		logarithm_table[1575] = 14'b0000011_1010000;
		logarithm_table[1576] = 14'b0000011_1010000;
		logarithm_table[1577] = 14'b0000011_1010000;
		logarithm_table[1578] = 14'b0000011_1010000;
		logarithm_table[1579] = 14'b0000011_1010000;
		logarithm_table[1580] = 14'b0000011_1010000;
		logarithm_table[1581] = 14'b0000011_1010000;
		logarithm_table[1582] = 14'b0000011_1010000;
		logarithm_table[1583] = 14'b0000011_1010000;
		logarithm_table[1584] = 14'b0000011_1010001;
		logarithm_table[1585] = 14'b0000011_1010001;
		logarithm_table[1586] = 14'b0000011_1010001;
		logarithm_table[1587] = 14'b0000011_1010001;
		logarithm_table[1588] = 14'b0000011_1010001;
		logarithm_table[1589] = 14'b0000011_1010001;
		logarithm_table[1590] = 14'b0000011_1010001;
		logarithm_table[1591] = 14'b0000011_1010001;
		logarithm_table[1592] = 14'b0000011_1010001;
		logarithm_table[1593] = 14'b0000011_1010010;
		logarithm_table[1594] = 14'b0000011_1010010;
		logarithm_table[1595] = 14'b0000011_1010010;
		logarithm_table[1596] = 14'b0000011_1010010;
		logarithm_table[1597] = 14'b0000011_1010010;
		logarithm_table[1598] = 14'b0000011_1010010;
		logarithm_table[1599] = 14'b0000011_1010010;
		logarithm_table[1600] = 14'b0000011_1010010;
		logarithm_table[1601] = 14'b0000011_1010011;
		logarithm_table[1602] = 14'b0000011_1010011;
		logarithm_table[1603] = 14'b0000011_1010011;
		logarithm_table[1604] = 14'b0000011_1010011;
		logarithm_table[1605] = 14'b0000011_1010011;
		logarithm_table[1606] = 14'b0000011_1010011;
		logarithm_table[1607] = 14'b0000011_1010011;
		logarithm_table[1608] = 14'b0000011_1010011;
		logarithm_table[1609] = 14'b0000011_1010011;
		logarithm_table[1610] = 14'b0000011_1010100;
		logarithm_table[1611] = 14'b0000011_1010100;
		logarithm_table[1612] = 14'b0000011_1010100;
		logarithm_table[1613] = 14'b0000011_1010100;
		logarithm_table[1614] = 14'b0000011_1010100;
		logarithm_table[1615] = 14'b0000011_1010100;
		logarithm_table[1616] = 14'b0000011_1010100;
		logarithm_table[1617] = 14'b0000011_1010100;
		logarithm_table[1618] = 14'b0000011_1010100;
		logarithm_table[1619] = 14'b0000011_1010101;
		logarithm_table[1620] = 14'b0000011_1010101;
		logarithm_table[1621] = 14'b0000011_1010101;
		logarithm_table[1622] = 14'b0000011_1010101;
		logarithm_table[1623] = 14'b0000011_1010101;
		logarithm_table[1624] = 14'b0000011_1010101;
		logarithm_table[1625] = 14'b0000011_1010101;
		logarithm_table[1626] = 14'b0000011_1010101;
		logarithm_table[1627] = 14'b0000011_1010110;
		logarithm_table[1628] = 14'b0000011_1010110;
		logarithm_table[1629] = 14'b0000011_1010110;
		logarithm_table[1630] = 14'b0000011_1010110;
		logarithm_table[1631] = 14'b0000011_1010110;
		logarithm_table[1632] = 14'b0000011_1010110;
		logarithm_table[1633] = 14'b0000011_1010110;
		logarithm_table[1634] = 14'b0000011_1010110;
		logarithm_table[1635] = 14'b0000011_1010110;
		logarithm_table[1636] = 14'b0000011_1010111;
		logarithm_table[1637] = 14'b0000011_1010111;
		logarithm_table[1638] = 14'b0000011_1010111;
		logarithm_table[1639] = 14'b0000011_1010111;
		logarithm_table[1640] = 14'b0000011_1010111;
		logarithm_table[1641] = 14'b0000011_1010111;
		logarithm_table[1642] = 14'b0000011_1010111;
		logarithm_table[1643] = 14'b0000011_1010111;
		logarithm_table[1644] = 14'b0000011_1010111;
		logarithm_table[1645] = 14'b0000011_1011000;
		logarithm_table[1646] = 14'b0000011_1011000;
		logarithm_table[1647] = 14'b0000011_1011000;
		logarithm_table[1648] = 14'b0000011_1011000;
		logarithm_table[1649] = 14'b0000011_1011000;
		logarithm_table[1650] = 14'b0000011_1011000;
		logarithm_table[1651] = 14'b0000011_1011000;
		logarithm_table[1652] = 14'b0000011_1011000;
		logarithm_table[1653] = 14'b0000011_1011000;
		logarithm_table[1654] = 14'b0000011_1011001;
		logarithm_table[1655] = 14'b0000011_1011001;
		logarithm_table[1656] = 14'b0000011_1011001;
		logarithm_table[1657] = 14'b0000011_1011001;
		logarithm_table[1658] = 14'b0000011_1011001;
		logarithm_table[1659] = 14'b0000011_1011001;
		logarithm_table[1660] = 14'b0000011_1011001;
		logarithm_table[1661] = 14'b0000011_1011001;
		logarithm_table[1662] = 14'b0000011_1011001;
		logarithm_table[1663] = 14'b0000011_1011010;
		logarithm_table[1664] = 14'b0000011_1011010;
		logarithm_table[1665] = 14'b0000011_1011010;
		logarithm_table[1666] = 14'b0000011_1011010;
		logarithm_table[1667] = 14'b0000011_1011010;
		logarithm_table[1668] = 14'b0000011_1011010;
		logarithm_table[1669] = 14'b0000011_1011010;
		logarithm_table[1670] = 14'b0000011_1011010;
		logarithm_table[1671] = 14'b0000011_1011010;
		logarithm_table[1672] = 14'b0000011_1011011;
		logarithm_table[1673] = 14'b0000011_1011011;
		logarithm_table[1674] = 14'b0000011_1011011;
		logarithm_table[1675] = 14'b0000011_1011011;
		logarithm_table[1676] = 14'b0000011_1011011;
		logarithm_table[1677] = 14'b0000011_1011011;
		logarithm_table[1678] = 14'b0000011_1011011;
		logarithm_table[1679] = 14'b0000011_1011011;
		logarithm_table[1680] = 14'b0000011_1011011;
		logarithm_table[1681] = 14'b0000011_1011100;
		logarithm_table[1682] = 14'b0000011_1011100;
		logarithm_table[1683] = 14'b0000011_1011100;
		logarithm_table[1684] = 14'b0000011_1011100;
		logarithm_table[1685] = 14'b0000011_1011100;
		logarithm_table[1686] = 14'b0000011_1011100;
		logarithm_table[1687] = 14'b0000011_1011100;
		logarithm_table[1688] = 14'b0000011_1011100;
		logarithm_table[1689] = 14'b0000011_1011100;
		logarithm_table[1690] = 14'b0000011_1011101;
		logarithm_table[1691] = 14'b0000011_1011101;
		logarithm_table[1692] = 14'b0000011_1011101;
		logarithm_table[1693] = 14'b0000011_1011101;
		logarithm_table[1694] = 14'b0000011_1011101;
		logarithm_table[1695] = 14'b0000011_1011101;
		logarithm_table[1696] = 14'b0000011_1011101;
		logarithm_table[1697] = 14'b0000011_1011101;
		logarithm_table[1698] = 14'b0000011_1011101;
		logarithm_table[1699] = 14'b0000011_1011110;
		logarithm_table[1700] = 14'b0000011_1011110;
		logarithm_table[1701] = 14'b0000011_1011110;
		logarithm_table[1702] = 14'b0000011_1011110;
		logarithm_table[1703] = 14'b0000011_1011110;
		logarithm_table[1704] = 14'b0000011_1011110;
		logarithm_table[1705] = 14'b0000011_1011110;
		logarithm_table[1706] = 14'b0000011_1011110;
		logarithm_table[1707] = 14'b0000011_1011110;
		logarithm_table[1708] = 14'b0000011_1011110;
		logarithm_table[1709] = 14'b0000011_1011111;
		logarithm_table[1710] = 14'b0000011_1011111;
		logarithm_table[1711] = 14'b0000011_1011111;
		logarithm_table[1712] = 14'b0000011_1011111;
		logarithm_table[1713] = 14'b0000011_1011111;
		logarithm_table[1714] = 14'b0000011_1011111;
		logarithm_table[1715] = 14'b0000011_1011111;
		logarithm_table[1716] = 14'b0000011_1011111;
		logarithm_table[1717] = 14'b0000011_1011111;
		logarithm_table[1718] = 14'b0000011_1100000;
		logarithm_table[1719] = 14'b0000011_1100000;
		logarithm_table[1720] = 14'b0000011_1100000;
		logarithm_table[1721] = 14'b0000011_1100000;
		logarithm_table[1722] = 14'b0000011_1100000;
		logarithm_table[1723] = 14'b0000011_1100000;
		logarithm_table[1724] = 14'b0000011_1100000;
		logarithm_table[1725] = 14'b0000011_1100000;
		logarithm_table[1726] = 14'b0000011_1100000;
		logarithm_table[1727] = 14'b0000011_1100001;
		logarithm_table[1728] = 14'b0000011_1100001;
		logarithm_table[1729] = 14'b0000011_1100001;
		logarithm_table[1730] = 14'b0000011_1100001;
		logarithm_table[1731] = 14'b0000011_1100001;
		logarithm_table[1732] = 14'b0000011_1100001;
		logarithm_table[1733] = 14'b0000011_1100001;
		logarithm_table[1734] = 14'b0000011_1100001;
		logarithm_table[1735] = 14'b0000011_1100001;
		logarithm_table[1736] = 14'b0000011_1100001;
		logarithm_table[1737] = 14'b0000011_1100010;
		logarithm_table[1738] = 14'b0000011_1100010;
		logarithm_table[1739] = 14'b0000011_1100010;
		logarithm_table[1740] = 14'b0000011_1100010;
		logarithm_table[1741] = 14'b0000011_1100010;
		logarithm_table[1742] = 14'b0000011_1100010;
		logarithm_table[1743] = 14'b0000011_1100010;
		logarithm_table[1744] = 14'b0000011_1100010;
		logarithm_table[1745] = 14'b0000011_1100010;
		logarithm_table[1746] = 14'b0000011_1100011;
		logarithm_table[1747] = 14'b0000011_1100011;
		logarithm_table[1748] = 14'b0000011_1100011;
		logarithm_table[1749] = 14'b0000011_1100011;
		logarithm_table[1750] = 14'b0000011_1100011;
		logarithm_table[1751] = 14'b0000011_1100011;
		logarithm_table[1752] = 14'b0000011_1100011;
		logarithm_table[1753] = 14'b0000011_1100011;
		logarithm_table[1754] = 14'b0000011_1100011;
		logarithm_table[1755] = 14'b0000011_1100011;
		logarithm_table[1756] = 14'b0000011_1100100;
		logarithm_table[1757] = 14'b0000011_1100100;
		logarithm_table[1758] = 14'b0000011_1100100;
		logarithm_table[1759] = 14'b0000011_1100100;
		logarithm_table[1760] = 14'b0000011_1100100;
		logarithm_table[1761] = 14'b0000011_1100100;
		logarithm_table[1762] = 14'b0000011_1100100;
		logarithm_table[1763] = 14'b0000011_1100100;
		logarithm_table[1764] = 14'b0000011_1100100;
		logarithm_table[1765] = 14'b0000011_1100101;
		logarithm_table[1766] = 14'b0000011_1100101;
		logarithm_table[1767] = 14'b0000011_1100101;
		logarithm_table[1768] = 14'b0000011_1100101;
		logarithm_table[1769] = 14'b0000011_1100101;
		logarithm_table[1770] = 14'b0000011_1100101;
		logarithm_table[1771] = 14'b0000011_1100101;
		logarithm_table[1772] = 14'b0000011_1100101;
		logarithm_table[1773] = 14'b0000011_1100101;
		logarithm_table[1774] = 14'b0000011_1100101;
		logarithm_table[1775] = 14'b0000011_1100110;
		logarithm_table[1776] = 14'b0000011_1100110;
		logarithm_table[1777] = 14'b0000011_1100110;
		logarithm_table[1778] = 14'b0000011_1100110;
		logarithm_table[1779] = 14'b0000011_1100110;
		logarithm_table[1780] = 14'b0000011_1100110;
		logarithm_table[1781] = 14'b0000011_1100110;
		logarithm_table[1782] = 14'b0000011_1100110;
		logarithm_table[1783] = 14'b0000011_1100110;
		logarithm_table[1784] = 14'b0000011_1100111;
		logarithm_table[1785] = 14'b0000011_1100111;
		logarithm_table[1786] = 14'b0000011_1100111;
		logarithm_table[1787] = 14'b0000011_1100111;
		logarithm_table[1788] = 14'b0000011_1100111;
		logarithm_table[1789] = 14'b0000011_1100111;
		logarithm_table[1790] = 14'b0000011_1100111;
		logarithm_table[1791] = 14'b0000011_1100111;
		logarithm_table[1792] = 14'b0000011_1100111;
		logarithm_table[1793] = 14'b0000011_1100111;
		logarithm_table[1794] = 14'b0000011_1101000;
		logarithm_table[1795] = 14'b0000011_1101000;
		logarithm_table[1796] = 14'b0000011_1101000;
		logarithm_table[1797] = 14'b0000011_1101000;
		logarithm_table[1798] = 14'b0000011_1101000;
		logarithm_table[1799] = 14'b0000011_1101000;
		logarithm_table[1800] = 14'b0000011_1101000;
		logarithm_table[1801] = 14'b0000011_1101000;
		logarithm_table[1802] = 14'b0000011_1101000;
		logarithm_table[1803] = 14'b0000011_1101000;
		logarithm_table[1804] = 14'b0000011_1101001;
		logarithm_table[1805] = 14'b0000011_1101001;
		logarithm_table[1806] = 14'b0000011_1101001;
		logarithm_table[1807] = 14'b0000011_1101001;
		logarithm_table[1808] = 14'b0000011_1101001;
		logarithm_table[1809] = 14'b0000011_1101001;
		logarithm_table[1810] = 14'b0000011_1101001;
		logarithm_table[1811] = 14'b0000011_1101001;
		logarithm_table[1812] = 14'b0000011_1101001;
		logarithm_table[1813] = 14'b0000011_1101001;
		logarithm_table[1814] = 14'b0000011_1101010;
		logarithm_table[1815] = 14'b0000011_1101010;
		logarithm_table[1816] = 14'b0000011_1101010;
		logarithm_table[1817] = 14'b0000011_1101010;
		logarithm_table[1818] = 14'b0000011_1101010;
		logarithm_table[1819] = 14'b0000011_1101010;
		logarithm_table[1820] = 14'b0000011_1101010;
		logarithm_table[1821] = 14'b0000011_1101010;
		logarithm_table[1822] = 14'b0000011_1101010;
		logarithm_table[1823] = 14'b0000011_1101011;
		logarithm_table[1824] = 14'b0000011_1101011;
		logarithm_table[1825] = 14'b0000011_1101011;
		logarithm_table[1826] = 14'b0000011_1101011;
		logarithm_table[1827] = 14'b0000011_1101011;
		logarithm_table[1828] = 14'b0000011_1101011;
		logarithm_table[1829] = 14'b0000011_1101011;
		logarithm_table[1830] = 14'b0000011_1101011;
		logarithm_table[1831] = 14'b0000011_1101011;
		logarithm_table[1832] = 14'b0000011_1101011;
		logarithm_table[1833] = 14'b0000011_1101100;
		logarithm_table[1834] = 14'b0000011_1101100;
		logarithm_table[1835] = 14'b0000011_1101100;
		logarithm_table[1836] = 14'b0000011_1101100;
		logarithm_table[1837] = 14'b0000011_1101100;
		logarithm_table[1838] = 14'b0000011_1101100;
		logarithm_table[1839] = 14'b0000011_1101100;
		logarithm_table[1840] = 14'b0000011_1101100;
		logarithm_table[1841] = 14'b0000011_1101100;
		logarithm_table[1842] = 14'b0000011_1101100;
		logarithm_table[1843] = 14'b0000011_1101101;
		logarithm_table[1844] = 14'b0000011_1101101;
		logarithm_table[1845] = 14'b0000011_1101101;
		logarithm_table[1846] = 14'b0000011_1101101;
		logarithm_table[1847] = 14'b0000011_1101101;
		logarithm_table[1848] = 14'b0000011_1101101;
		logarithm_table[1849] = 14'b0000011_1101101;
		logarithm_table[1850] = 14'b0000011_1101101;
		logarithm_table[1851] = 14'b0000011_1101101;
		logarithm_table[1852] = 14'b0000011_1101101;
		logarithm_table[1853] = 14'b0000011_1101110;
		logarithm_table[1854] = 14'b0000011_1101110;
		logarithm_table[1855] = 14'b0000011_1101110;
		logarithm_table[1856] = 14'b0000011_1101110;
		logarithm_table[1857] = 14'b0000011_1101110;
		logarithm_table[1858] = 14'b0000011_1101110;
		logarithm_table[1859] = 14'b0000011_1101110;
		logarithm_table[1860] = 14'b0000011_1101110;
		logarithm_table[1861] = 14'b0000011_1101110;
		logarithm_table[1862] = 14'b0000011_1101110;
		logarithm_table[1863] = 14'b0000011_1101111;
		logarithm_table[1864] = 14'b0000011_1101111;
		logarithm_table[1865] = 14'b0000011_1101111;
		logarithm_table[1866] = 14'b0000011_1101111;
		logarithm_table[1867] = 14'b0000011_1101111;
		logarithm_table[1868] = 14'b0000011_1101111;
		logarithm_table[1869] = 14'b0000011_1101111;
		logarithm_table[1870] = 14'b0000011_1101111;
		logarithm_table[1871] = 14'b0000011_1101111;
		logarithm_table[1872] = 14'b0000011_1101111;
		logarithm_table[1873] = 14'b0000011_1110000;
		logarithm_table[1874] = 14'b0000011_1110000;
		logarithm_table[1875] = 14'b0000011_1110000;
		logarithm_table[1876] = 14'b0000011_1110000;
		logarithm_table[1877] = 14'b0000011_1110000;
		logarithm_table[1878] = 14'b0000011_1110000;
		logarithm_table[1879] = 14'b0000011_1110000;
		logarithm_table[1880] = 14'b0000011_1110000;
		logarithm_table[1881] = 14'b0000011_1110000;
		logarithm_table[1882] = 14'b0000011_1110000;
		logarithm_table[1883] = 14'b0000011_1110000;
		logarithm_table[1884] = 14'b0000011_1110001;
		logarithm_table[1885] = 14'b0000011_1110001;
		logarithm_table[1886] = 14'b0000011_1110001;
		logarithm_table[1887] = 14'b0000011_1110001;
		logarithm_table[1888] = 14'b0000011_1110001;
		logarithm_table[1889] = 14'b0000011_1110001;
		logarithm_table[1890] = 14'b0000011_1110001;
		logarithm_table[1891] = 14'b0000011_1110001;
		logarithm_table[1892] = 14'b0000011_1110001;
		logarithm_table[1893] = 14'b0000011_1110001;
		logarithm_table[1894] = 14'b0000011_1110010;
		logarithm_table[1895] = 14'b0000011_1110010;
		logarithm_table[1896] = 14'b0000011_1110010;
		logarithm_table[1897] = 14'b0000011_1110010;
		logarithm_table[1898] = 14'b0000011_1110010;
		logarithm_table[1899] = 14'b0000011_1110010;
		logarithm_table[1900] = 14'b0000011_1110010;
		logarithm_table[1901] = 14'b0000011_1110010;
		logarithm_table[1902] = 14'b0000011_1110010;
		logarithm_table[1903] = 14'b0000011_1110010;
		logarithm_table[1904] = 14'b0000011_1110011;
		logarithm_table[1905] = 14'b0000011_1110011;
		logarithm_table[1906] = 14'b0000011_1110011;
		logarithm_table[1907] = 14'b0000011_1110011;
		logarithm_table[1908] = 14'b0000011_1110011;
		logarithm_table[1909] = 14'b0000011_1110011;
		logarithm_table[1910] = 14'b0000011_1110011;
		logarithm_table[1911] = 14'b0000011_1110011;
		logarithm_table[1912] = 14'b0000011_1110011;
		logarithm_table[1913] = 14'b0000011_1110011;
		logarithm_table[1914] = 14'b0000011_1110100;
		logarithm_table[1915] = 14'b0000011_1110100;
		logarithm_table[1916] = 14'b0000011_1110100;
		logarithm_table[1917] = 14'b0000011_1110100;
		logarithm_table[1918] = 14'b0000011_1110100;
		logarithm_table[1919] = 14'b0000011_1110100;
		logarithm_table[1920] = 14'b0000011_1110100;
		logarithm_table[1921] = 14'b0000011_1110100;
		logarithm_table[1922] = 14'b0000011_1110100;
		logarithm_table[1923] = 14'b0000011_1110100;
		logarithm_table[1924] = 14'b0000011_1110100;
		logarithm_table[1925] = 14'b0000011_1110101;
		logarithm_table[1926] = 14'b0000011_1110101;
		logarithm_table[1927] = 14'b0000011_1110101;
		logarithm_table[1928] = 14'b0000011_1110101;
		logarithm_table[1929] = 14'b0000011_1110101;
		logarithm_table[1930] = 14'b0000011_1110101;
		logarithm_table[1931] = 14'b0000011_1110101;
		logarithm_table[1932] = 14'b0000011_1110101;
		logarithm_table[1933] = 14'b0000011_1110101;
		logarithm_table[1934] = 14'b0000011_1110101;
		logarithm_table[1935] = 14'b0000011_1110110;
		logarithm_table[1936] = 14'b0000011_1110110;
		logarithm_table[1937] = 14'b0000011_1110110;
		logarithm_table[1938] = 14'b0000011_1110110;
		logarithm_table[1939] = 14'b0000011_1110110;
		logarithm_table[1940] = 14'b0000011_1110110;
		logarithm_table[1941] = 14'b0000011_1110110;
		logarithm_table[1942] = 14'b0000011_1110110;
		logarithm_table[1943] = 14'b0000011_1110110;
		logarithm_table[1944] = 14'b0000011_1110110;
		logarithm_table[1945] = 14'b0000011_1110110;
		logarithm_table[1946] = 14'b0000011_1110111;
		logarithm_table[1947] = 14'b0000011_1110111;
		logarithm_table[1948] = 14'b0000011_1110111;
		logarithm_table[1949] = 14'b0000011_1110111;
		logarithm_table[1950] = 14'b0000011_1110111;
		logarithm_table[1951] = 14'b0000011_1110111;
		logarithm_table[1952] = 14'b0000011_1110111;
		logarithm_table[1953] = 14'b0000011_1110111;
		logarithm_table[1954] = 14'b0000011_1110111;
		logarithm_table[1955] = 14'b0000011_1110111;
		logarithm_table[1956] = 14'b0000011_1111000;
		logarithm_table[1957] = 14'b0000011_1111000;
		logarithm_table[1958] = 14'b0000011_1111000;
		logarithm_table[1959] = 14'b0000011_1111000;
		logarithm_table[1960] = 14'b0000011_1111000;
		logarithm_table[1961] = 14'b0000011_1111000;
		logarithm_table[1962] = 14'b0000011_1111000;
		logarithm_table[1963] = 14'b0000011_1111000;
		logarithm_table[1964] = 14'b0000011_1111000;
		logarithm_table[1965] = 14'b0000011_1111000;
		logarithm_table[1966] = 14'b0000011_1111000;
		logarithm_table[1967] = 14'b0000011_1111001;
		logarithm_table[1968] = 14'b0000011_1111001;
		logarithm_table[1969] = 14'b0000011_1111001;
		logarithm_table[1970] = 14'b0000011_1111001;
		logarithm_table[1971] = 14'b0000011_1111001;
		logarithm_table[1972] = 14'b0000011_1111001;
		logarithm_table[1973] = 14'b0000011_1111001;
		logarithm_table[1974] = 14'b0000011_1111001;
		logarithm_table[1975] = 14'b0000011_1111001;
		logarithm_table[1976] = 14'b0000011_1111001;
		logarithm_table[1977] = 14'b0000011_1111001;
		logarithm_table[1978] = 14'b0000011_1111010;
		logarithm_table[1979] = 14'b0000011_1111010;
		logarithm_table[1980] = 14'b0000011_1111010;
		logarithm_table[1981] = 14'b0000011_1111010;
		logarithm_table[1982] = 14'b0000011_1111010;
		logarithm_table[1983] = 14'b0000011_1111010;
		logarithm_table[1984] = 14'b0000011_1111010;
		logarithm_table[1985] = 14'b0000011_1111010;
		logarithm_table[1986] = 14'b0000011_1111010;
		logarithm_table[1987] = 14'b0000011_1111010;
		logarithm_table[1988] = 14'b0000011_1111011;
		logarithm_table[1989] = 14'b0000011_1111011;
		logarithm_table[1990] = 14'b0000011_1111011;
		logarithm_table[1991] = 14'b0000011_1111011;
		logarithm_table[1992] = 14'b0000011_1111011;
		logarithm_table[1993] = 14'b0000011_1111011;
		logarithm_table[1994] = 14'b0000011_1111011;
		logarithm_table[1995] = 14'b0000011_1111011;
		logarithm_table[1996] = 14'b0000011_1111011;
		logarithm_table[1997] = 14'b0000011_1111011;
		logarithm_table[1998] = 14'b0000011_1111011;
		logarithm_table[1999] = 14'b0000011_1111100;
		logarithm_table[2000] = 14'b0000011_1111100;
		logarithm_table[2001] = 14'b0000011_1111100;
		logarithm_table[2002] = 14'b0000011_1111100;
		logarithm_table[2003] = 14'b0000011_1111100;
		logarithm_table[2004] = 14'b0000011_1111100;
		logarithm_table[2005] = 14'b0000011_1111100;
		logarithm_table[2006] = 14'b0000011_1111100;
		logarithm_table[2007] = 14'b0000011_1111100;
		logarithm_table[2008] = 14'b0000011_1111100;
		logarithm_table[2009] = 14'b0000011_1111100;
		logarithm_table[2010] = 14'b0000011_1111101;
		logarithm_table[2011] = 14'b0000011_1111101;
		logarithm_table[2012] = 14'b0000011_1111101;
		logarithm_table[2013] = 14'b0000011_1111101;
		logarithm_table[2014] = 14'b0000011_1111101;
		logarithm_table[2015] = 14'b0000011_1111101;
		logarithm_table[2016] = 14'b0000011_1111101;
		logarithm_table[2017] = 14'b0000011_1111101;
		logarithm_table[2018] = 14'b0000011_1111101;
		logarithm_table[2019] = 14'b0000011_1111101;
		logarithm_table[2020] = 14'b0000011_1111101;
		logarithm_table[2021] = 14'b0000011_1111110;
		logarithm_table[2022] = 14'b0000011_1111110;
		logarithm_table[2023] = 14'b0000011_1111110;
		logarithm_table[2024] = 14'b0000011_1111110;
		logarithm_table[2025] = 14'b0000011_1111110;
		logarithm_table[2026] = 14'b0000011_1111110;
		logarithm_table[2027] = 14'b0000011_1111110;
		logarithm_table[2028] = 14'b0000011_1111110;
		logarithm_table[2029] = 14'b0000011_1111110;
		logarithm_table[2030] = 14'b0000011_1111110;
		logarithm_table[2031] = 14'b0000011_1111110;
		logarithm_table[2032] = 14'b0000011_1111111;
		logarithm_table[2033] = 14'b0000011_1111111;
		logarithm_table[2034] = 14'b0000011_1111111;
		logarithm_table[2035] = 14'b0000011_1111111;
		logarithm_table[2036] = 14'b0000011_1111111;
		logarithm_table[2037] = 14'b0000011_1111111;
		logarithm_table[2038] = 14'b0000011_1111111;
		logarithm_table[2039] = 14'b0000011_1111111;
		logarithm_table[2040] = 14'b0000011_1111111;
		logarithm_table[2041] = 14'b0000011_1111111;
		logarithm_table[2042] = 14'b0000011_1111111;
		logarithm_table[2043] = 14'b0000100_0000000;
		logarithm_table[2044] = 14'b0000100_0000000;
		logarithm_table[2045] = 14'b0000100_0000000;
		logarithm_table[2046] = 14'b0000100_0000000;
		logarithm_table[2047] = 14'b0000100_0000000;
		logarithm_table[2048] = 14'b0000100_0000000;
		logarithm_table[2049] = 14'b0000100_0000000;
		logarithm_table[2050] = 14'b0000100_0000000;
		logarithm_table[2051] = 14'b0000100_0000000;
		logarithm_table[2052] = 14'b0000100_0000000;
		logarithm_table[2053] = 14'b0000100_0000000;
		logarithm_table[2054] = 14'b0000100_0000001;
		logarithm_table[2055] = 14'b0000100_0000001;
		logarithm_table[2056] = 14'b0000100_0000001;
		logarithm_table[2057] = 14'b0000100_0000001;
		logarithm_table[2058] = 14'b0000100_0000001;
		logarithm_table[2059] = 14'b0000100_0000001;
		logarithm_table[2060] = 14'b0000100_0000001;
		logarithm_table[2061] = 14'b0000100_0000001;
		logarithm_table[2062] = 14'b0000100_0000001;
		logarithm_table[2063] = 14'b0000100_0000001;
		logarithm_table[2064] = 14'b0000100_0000001;
		logarithm_table[2065] = 14'b0000100_0000010;
		logarithm_table[2066] = 14'b0000100_0000010;
		logarithm_table[2067] = 14'b0000100_0000010;
		logarithm_table[2068] = 14'b0000100_0000010;
		logarithm_table[2069] = 14'b0000100_0000010;
		logarithm_table[2070] = 14'b0000100_0000010;
		logarithm_table[2071] = 14'b0000100_0000010;
		logarithm_table[2072] = 14'b0000100_0000010;
		logarithm_table[2073] = 14'b0000100_0000010;
		logarithm_table[2074] = 14'b0000100_0000010;
		logarithm_table[2075] = 14'b0000100_0000010;
		logarithm_table[2076] = 14'b0000100_0000011;
		logarithm_table[2077] = 14'b0000100_0000011;
		logarithm_table[2078] = 14'b0000100_0000011;
		logarithm_table[2079] = 14'b0000100_0000011;
		logarithm_table[2080] = 14'b0000100_0000011;
		logarithm_table[2081] = 14'b0000100_0000011;
		logarithm_table[2082] = 14'b0000100_0000011;
		logarithm_table[2083] = 14'b0000100_0000011;
		logarithm_table[2084] = 14'b0000100_0000011;
		logarithm_table[2085] = 14'b0000100_0000011;
		logarithm_table[2086] = 14'b0000100_0000011;
		logarithm_table[2087] = 14'b0000100_0000011;
		logarithm_table[2088] = 14'b0000100_0000100;
		logarithm_table[2089] = 14'b0000100_0000100;
		logarithm_table[2090] = 14'b0000100_0000100;
		logarithm_table[2091] = 14'b0000100_0000100;
		logarithm_table[2092] = 14'b0000100_0000100;
		logarithm_table[2093] = 14'b0000100_0000100;
		logarithm_table[2094] = 14'b0000100_0000100;
		logarithm_table[2095] = 14'b0000100_0000100;
		logarithm_table[2096] = 14'b0000100_0000100;
		logarithm_table[2097] = 14'b0000100_0000100;
		logarithm_table[2098] = 14'b0000100_0000100;
		logarithm_table[2099] = 14'b0000100_0000101;
		logarithm_table[2100] = 14'b0000100_0000101;
		logarithm_table[2101] = 14'b0000100_0000101;
		logarithm_table[2102] = 14'b0000100_0000101;
		logarithm_table[2103] = 14'b0000100_0000101;
		logarithm_table[2104] = 14'b0000100_0000101;
		logarithm_table[2105] = 14'b0000100_0000101;
		logarithm_table[2106] = 14'b0000100_0000101;
		logarithm_table[2107] = 14'b0000100_0000101;
		logarithm_table[2108] = 14'b0000100_0000101;
		logarithm_table[2109] = 14'b0000100_0000101;
		logarithm_table[2110] = 14'b0000100_0000110;
		logarithm_table[2111] = 14'b0000100_0000110;
		logarithm_table[2112] = 14'b0000100_0000110;
		logarithm_table[2113] = 14'b0000100_0000110;
		logarithm_table[2114] = 14'b0000100_0000110;
		logarithm_table[2115] = 14'b0000100_0000110;
		logarithm_table[2116] = 14'b0000100_0000110;
		logarithm_table[2117] = 14'b0000100_0000110;
		logarithm_table[2118] = 14'b0000100_0000110;
		logarithm_table[2119] = 14'b0000100_0000110;
		logarithm_table[2120] = 14'b0000100_0000110;
		logarithm_table[2121] = 14'b0000100_0000110;
		logarithm_table[2122] = 14'b0000100_0000111;
		logarithm_table[2123] = 14'b0000100_0000111;
		logarithm_table[2124] = 14'b0000100_0000111;
		logarithm_table[2125] = 14'b0000100_0000111;
		logarithm_table[2126] = 14'b0000100_0000111;
		logarithm_table[2127] = 14'b0000100_0000111;
		logarithm_table[2128] = 14'b0000100_0000111;
		logarithm_table[2129] = 14'b0000100_0000111;
		logarithm_table[2130] = 14'b0000100_0000111;
		logarithm_table[2131] = 14'b0000100_0000111;
		logarithm_table[2132] = 14'b0000100_0000111;
		logarithm_table[2133] = 14'b0000100_0001000;
		logarithm_table[2134] = 14'b0000100_0001000;
		logarithm_table[2135] = 14'b0000100_0001000;
		logarithm_table[2136] = 14'b0000100_0001000;
		logarithm_table[2137] = 14'b0000100_0001000;
		logarithm_table[2138] = 14'b0000100_0001000;
		logarithm_table[2139] = 14'b0000100_0001000;
		logarithm_table[2140] = 14'b0000100_0001000;
		logarithm_table[2141] = 14'b0000100_0001000;
		logarithm_table[2142] = 14'b0000100_0001000;
		logarithm_table[2143] = 14'b0000100_0001000;
		logarithm_table[2144] = 14'b0000100_0001000;
		logarithm_table[2145] = 14'b0000100_0001001;
		logarithm_table[2146] = 14'b0000100_0001001;
		logarithm_table[2147] = 14'b0000100_0001001;
		logarithm_table[2148] = 14'b0000100_0001001;
		logarithm_table[2149] = 14'b0000100_0001001;
		logarithm_table[2150] = 14'b0000100_0001001;
		logarithm_table[2151] = 14'b0000100_0001001;
		logarithm_table[2152] = 14'b0000100_0001001;
		logarithm_table[2153] = 14'b0000100_0001001;
		logarithm_table[2154] = 14'b0000100_0001001;
		logarithm_table[2155] = 14'b0000100_0001001;
		logarithm_table[2156] = 14'b0000100_0001001;
		logarithm_table[2157] = 14'b0000100_0001010;
		logarithm_table[2158] = 14'b0000100_0001010;
		logarithm_table[2159] = 14'b0000100_0001010;
		logarithm_table[2160] = 14'b0000100_0001010;
		logarithm_table[2161] = 14'b0000100_0001010;
		logarithm_table[2162] = 14'b0000100_0001010;
		logarithm_table[2163] = 14'b0000100_0001010;
		logarithm_table[2164] = 14'b0000100_0001010;
		logarithm_table[2165] = 14'b0000100_0001010;
		logarithm_table[2166] = 14'b0000100_0001010;
		logarithm_table[2167] = 14'b0000100_0001010;
		logarithm_table[2168] = 14'b0000100_0001011;
		logarithm_table[2169] = 14'b0000100_0001011;
		logarithm_table[2170] = 14'b0000100_0001011;
		logarithm_table[2171] = 14'b0000100_0001011;
		logarithm_table[2172] = 14'b0000100_0001011;
		logarithm_table[2173] = 14'b0000100_0001011;
		logarithm_table[2174] = 14'b0000100_0001011;
		logarithm_table[2175] = 14'b0000100_0001011;
		logarithm_table[2176] = 14'b0000100_0001011;
		logarithm_table[2177] = 14'b0000100_0001011;
		logarithm_table[2178] = 14'b0000100_0001011;
		logarithm_table[2179] = 14'b0000100_0001011;
		logarithm_table[2180] = 14'b0000100_0001100;
		logarithm_table[2181] = 14'b0000100_0001100;
		logarithm_table[2182] = 14'b0000100_0001100;
		logarithm_table[2183] = 14'b0000100_0001100;
		logarithm_table[2184] = 14'b0000100_0001100;
		logarithm_table[2185] = 14'b0000100_0001100;
		logarithm_table[2186] = 14'b0000100_0001100;
		logarithm_table[2187] = 14'b0000100_0001100;
		logarithm_table[2188] = 14'b0000100_0001100;
		logarithm_table[2189] = 14'b0000100_0001100;
		logarithm_table[2190] = 14'b0000100_0001100;
		logarithm_table[2191] = 14'b0000100_0001100;
		logarithm_table[2192] = 14'b0000100_0001101;
		logarithm_table[2193] = 14'b0000100_0001101;
		logarithm_table[2194] = 14'b0000100_0001101;
		logarithm_table[2195] = 14'b0000100_0001101;
		logarithm_table[2196] = 14'b0000100_0001101;
		logarithm_table[2197] = 14'b0000100_0001101;
		logarithm_table[2198] = 14'b0000100_0001101;
		logarithm_table[2199] = 14'b0000100_0001101;
		logarithm_table[2200] = 14'b0000100_0001101;
		logarithm_table[2201] = 14'b0000100_0001101;
		logarithm_table[2202] = 14'b0000100_0001101;
		logarithm_table[2203] = 14'b0000100_0001101;
		logarithm_table[2204] = 14'b0000100_0001110;
		logarithm_table[2205] = 14'b0000100_0001110;
		logarithm_table[2206] = 14'b0000100_0001110;
		logarithm_table[2207] = 14'b0000100_0001110;
		logarithm_table[2208] = 14'b0000100_0001110;
		logarithm_table[2209] = 14'b0000100_0001110;
		logarithm_table[2210] = 14'b0000100_0001110;
		logarithm_table[2211] = 14'b0000100_0001110;
		logarithm_table[2212] = 14'b0000100_0001110;
		logarithm_table[2213] = 14'b0000100_0001110;
		logarithm_table[2214] = 14'b0000100_0001110;
		logarithm_table[2215] = 14'b0000100_0001110;
		logarithm_table[2216] = 14'b0000100_0001111;
		logarithm_table[2217] = 14'b0000100_0001111;
		logarithm_table[2218] = 14'b0000100_0001111;
		logarithm_table[2219] = 14'b0000100_0001111;
		logarithm_table[2220] = 14'b0000100_0001111;
		logarithm_table[2221] = 14'b0000100_0001111;
		logarithm_table[2222] = 14'b0000100_0001111;
		logarithm_table[2223] = 14'b0000100_0001111;
		logarithm_table[2224] = 14'b0000100_0001111;
		logarithm_table[2225] = 14'b0000100_0001111;
		logarithm_table[2226] = 14'b0000100_0001111;
		logarithm_table[2227] = 14'b0000100_0001111;
		logarithm_table[2228] = 14'b0000100_0010000;
		logarithm_table[2229] = 14'b0000100_0010000;
		logarithm_table[2230] = 14'b0000100_0010000;
		logarithm_table[2231] = 14'b0000100_0010000;
		logarithm_table[2232] = 14'b0000100_0010000;
		logarithm_table[2233] = 14'b0000100_0010000;
		logarithm_table[2234] = 14'b0000100_0010000;
		logarithm_table[2235] = 14'b0000100_0010000;
		logarithm_table[2236] = 14'b0000100_0010000;
		logarithm_table[2237] = 14'b0000100_0010000;
		logarithm_table[2238] = 14'b0000100_0010000;
		logarithm_table[2239] = 14'b0000100_0010000;
		logarithm_table[2240] = 14'b0000100_0010001;
		logarithm_table[2241] = 14'b0000100_0010001;
		logarithm_table[2242] = 14'b0000100_0010001;
		logarithm_table[2243] = 14'b0000100_0010001;
		logarithm_table[2244] = 14'b0000100_0010001;
		logarithm_table[2245] = 14'b0000100_0010001;
		logarithm_table[2246] = 14'b0000100_0010001;
		logarithm_table[2247] = 14'b0000100_0010001;
		logarithm_table[2248] = 14'b0000100_0010001;
		logarithm_table[2249] = 14'b0000100_0010001;
		logarithm_table[2250] = 14'b0000100_0010001;
		logarithm_table[2251] = 14'b0000100_0010001;
		logarithm_table[2252] = 14'b0000100_0010010;
		logarithm_table[2253] = 14'b0000100_0010010;
		logarithm_table[2254] = 14'b0000100_0010010;
		logarithm_table[2255] = 14'b0000100_0010010;
		logarithm_table[2256] = 14'b0000100_0010010;
		logarithm_table[2257] = 14'b0000100_0010010;
		logarithm_table[2258] = 14'b0000100_0010010;
		logarithm_table[2259] = 14'b0000100_0010010;
		logarithm_table[2260] = 14'b0000100_0010010;
		logarithm_table[2261] = 14'b0000100_0010010;
		logarithm_table[2262] = 14'b0000100_0010010;
		logarithm_table[2263] = 14'b0000100_0010010;
		logarithm_table[2264] = 14'b0000100_0010011;
		logarithm_table[2265] = 14'b0000100_0010011;
		logarithm_table[2266] = 14'b0000100_0010011;
		logarithm_table[2267] = 14'b0000100_0010011;
		logarithm_table[2268] = 14'b0000100_0010011;
		logarithm_table[2269] = 14'b0000100_0010011;
		logarithm_table[2270] = 14'b0000100_0010011;
		logarithm_table[2271] = 14'b0000100_0010011;
		logarithm_table[2272] = 14'b0000100_0010011;
		logarithm_table[2273] = 14'b0000100_0010011;
		logarithm_table[2274] = 14'b0000100_0010011;
		logarithm_table[2275] = 14'b0000100_0010011;
		logarithm_table[2276] = 14'b0000100_0010011;
		logarithm_table[2277] = 14'b0000100_0010100;
		logarithm_table[2278] = 14'b0000100_0010100;
		logarithm_table[2279] = 14'b0000100_0010100;
		logarithm_table[2280] = 14'b0000100_0010100;
		logarithm_table[2281] = 14'b0000100_0010100;
		logarithm_table[2282] = 14'b0000100_0010100;
		logarithm_table[2283] = 14'b0000100_0010100;
		logarithm_table[2284] = 14'b0000100_0010100;
		logarithm_table[2285] = 14'b0000100_0010100;
		logarithm_table[2286] = 14'b0000100_0010100;
		logarithm_table[2287] = 14'b0000100_0010100;
		logarithm_table[2288] = 14'b0000100_0010100;
		logarithm_table[2289] = 14'b0000100_0010101;
		logarithm_table[2290] = 14'b0000100_0010101;
		logarithm_table[2291] = 14'b0000100_0010101;
		logarithm_table[2292] = 14'b0000100_0010101;
		logarithm_table[2293] = 14'b0000100_0010101;
		logarithm_table[2294] = 14'b0000100_0010101;
		logarithm_table[2295] = 14'b0000100_0010101;
		logarithm_table[2296] = 14'b0000100_0010101;
		logarithm_table[2297] = 14'b0000100_0010101;
		logarithm_table[2298] = 14'b0000100_0010101;
		logarithm_table[2299] = 14'b0000100_0010101;
		logarithm_table[2300] = 14'b0000100_0010101;
		logarithm_table[2301] = 14'b0000100_0010110;
		logarithm_table[2302] = 14'b0000100_0010110;
		logarithm_table[2303] = 14'b0000100_0010110;
		logarithm_table[2304] = 14'b0000100_0010110;
		logarithm_table[2305] = 14'b0000100_0010110;
		logarithm_table[2306] = 14'b0000100_0010110;
		logarithm_table[2307] = 14'b0000100_0010110;
		logarithm_table[2308] = 14'b0000100_0010110;
		logarithm_table[2309] = 14'b0000100_0010110;
		logarithm_table[2310] = 14'b0000100_0010110;
		logarithm_table[2311] = 14'b0000100_0010110;
		logarithm_table[2312] = 14'b0000100_0010110;
		logarithm_table[2313] = 14'b0000100_0010110;
		logarithm_table[2314] = 14'b0000100_0010111;
		logarithm_table[2315] = 14'b0000100_0010111;
		logarithm_table[2316] = 14'b0000100_0010111;
		logarithm_table[2317] = 14'b0000100_0010111;
		logarithm_table[2318] = 14'b0000100_0010111;
		logarithm_table[2319] = 14'b0000100_0010111;
		logarithm_table[2320] = 14'b0000100_0010111;
		logarithm_table[2321] = 14'b0000100_0010111;
		logarithm_table[2322] = 14'b0000100_0010111;
		logarithm_table[2323] = 14'b0000100_0010111;
		logarithm_table[2324] = 14'b0000100_0010111;
		logarithm_table[2325] = 14'b0000100_0010111;
		logarithm_table[2326] = 14'b0000100_0011000;
		logarithm_table[2327] = 14'b0000100_0011000;
		logarithm_table[2328] = 14'b0000100_0011000;
		logarithm_table[2329] = 14'b0000100_0011000;
		logarithm_table[2330] = 14'b0000100_0011000;
		logarithm_table[2331] = 14'b0000100_0011000;
		logarithm_table[2332] = 14'b0000100_0011000;
		logarithm_table[2333] = 14'b0000100_0011000;
		logarithm_table[2334] = 14'b0000100_0011000;
		logarithm_table[2335] = 14'b0000100_0011000;
		logarithm_table[2336] = 14'b0000100_0011000;
		logarithm_table[2337] = 14'b0000100_0011000;
		logarithm_table[2338] = 14'b0000100_0011000;
		logarithm_table[2339] = 14'b0000100_0011001;
		logarithm_table[2340] = 14'b0000100_0011001;
		logarithm_table[2341] = 14'b0000100_0011001;
		logarithm_table[2342] = 14'b0000100_0011001;
		logarithm_table[2343] = 14'b0000100_0011001;
		logarithm_table[2344] = 14'b0000100_0011001;
		logarithm_table[2345] = 14'b0000100_0011001;
		logarithm_table[2346] = 14'b0000100_0011001;
		logarithm_table[2347] = 14'b0000100_0011001;
		logarithm_table[2348] = 14'b0000100_0011001;
		logarithm_table[2349] = 14'b0000100_0011001;
		logarithm_table[2350] = 14'b0000100_0011001;
		logarithm_table[2351] = 14'b0000100_0011001;
		logarithm_table[2352] = 14'b0000100_0011010;
		logarithm_table[2353] = 14'b0000100_0011010;
		logarithm_table[2354] = 14'b0000100_0011010;
		logarithm_table[2355] = 14'b0000100_0011010;
		logarithm_table[2356] = 14'b0000100_0011010;
		logarithm_table[2357] = 14'b0000100_0011010;
		logarithm_table[2358] = 14'b0000100_0011010;
		logarithm_table[2359] = 14'b0000100_0011010;
		logarithm_table[2360] = 14'b0000100_0011010;
		logarithm_table[2361] = 14'b0000100_0011010;
		logarithm_table[2362] = 14'b0000100_0011010;
		logarithm_table[2363] = 14'b0000100_0011010;
		logarithm_table[2364] = 14'b0000100_0011010;
		logarithm_table[2365] = 14'b0000100_0011011;
		logarithm_table[2366] = 14'b0000100_0011011;
		logarithm_table[2367] = 14'b0000100_0011011;
		logarithm_table[2368] = 14'b0000100_0011011;
		logarithm_table[2369] = 14'b0000100_0011011;
		logarithm_table[2370] = 14'b0000100_0011011;
		logarithm_table[2371] = 14'b0000100_0011011;
		logarithm_table[2372] = 14'b0000100_0011011;
		logarithm_table[2373] = 14'b0000100_0011011;
		logarithm_table[2374] = 14'b0000100_0011011;
		logarithm_table[2375] = 14'b0000100_0011011;
		logarithm_table[2376] = 14'b0000100_0011011;
		logarithm_table[2377] = 14'b0000100_0011100;
		logarithm_table[2378] = 14'b0000100_0011100;
		logarithm_table[2379] = 14'b0000100_0011100;
		logarithm_table[2380] = 14'b0000100_0011100;
		logarithm_table[2381] = 14'b0000100_0011100;
		logarithm_table[2382] = 14'b0000100_0011100;
		logarithm_table[2383] = 14'b0000100_0011100;
		logarithm_table[2384] = 14'b0000100_0011100;
		logarithm_table[2385] = 14'b0000100_0011100;
		logarithm_table[2386] = 14'b0000100_0011100;
		logarithm_table[2387] = 14'b0000100_0011100;
		logarithm_table[2388] = 14'b0000100_0011100;
		logarithm_table[2389] = 14'b0000100_0011100;
		logarithm_table[2390] = 14'b0000100_0011101;
		logarithm_table[2391] = 14'b0000100_0011101;
		logarithm_table[2392] = 14'b0000100_0011101;
		logarithm_table[2393] = 14'b0000100_0011101;
		logarithm_table[2394] = 14'b0000100_0011101;
		logarithm_table[2395] = 14'b0000100_0011101;
		logarithm_table[2396] = 14'b0000100_0011101;
		logarithm_table[2397] = 14'b0000100_0011101;
		logarithm_table[2398] = 14'b0000100_0011101;
		logarithm_table[2399] = 14'b0000100_0011101;
		logarithm_table[2400] = 14'b0000100_0011101;
		logarithm_table[2401] = 14'b0000100_0011101;
		logarithm_table[2402] = 14'b0000100_0011101;
		logarithm_table[2403] = 14'b0000100_0011110;
		logarithm_table[2404] = 14'b0000100_0011110;
		logarithm_table[2405] = 14'b0000100_0011110;
		logarithm_table[2406] = 14'b0000100_0011110;
		logarithm_table[2407] = 14'b0000100_0011110;
		logarithm_table[2408] = 14'b0000100_0011110;
		logarithm_table[2409] = 14'b0000100_0011110;
		logarithm_table[2410] = 14'b0000100_0011110;
		logarithm_table[2411] = 14'b0000100_0011110;
		logarithm_table[2412] = 14'b0000100_0011110;
		logarithm_table[2413] = 14'b0000100_0011110;
		logarithm_table[2414] = 14'b0000100_0011110;
		logarithm_table[2415] = 14'b0000100_0011110;
		logarithm_table[2416] = 14'b0000100_0011111;
		logarithm_table[2417] = 14'b0000100_0011111;
		logarithm_table[2418] = 14'b0000100_0011111;
		logarithm_table[2419] = 14'b0000100_0011111;
		logarithm_table[2420] = 14'b0000100_0011111;
		logarithm_table[2421] = 14'b0000100_0011111;
		logarithm_table[2422] = 14'b0000100_0011111;
		logarithm_table[2423] = 14'b0000100_0011111;
		logarithm_table[2424] = 14'b0000100_0011111;
		logarithm_table[2425] = 14'b0000100_0011111;
		logarithm_table[2426] = 14'b0000100_0011111;
		logarithm_table[2427] = 14'b0000100_0011111;
		logarithm_table[2428] = 14'b0000100_0011111;
		logarithm_table[2429] = 14'b0000100_0100000;
		logarithm_table[2430] = 14'b0000100_0100000;
		logarithm_table[2431] = 14'b0000100_0100000;
		logarithm_table[2432] = 14'b0000100_0100000;
		logarithm_table[2433] = 14'b0000100_0100000;
		logarithm_table[2434] = 14'b0000100_0100000;
		logarithm_table[2435] = 14'b0000100_0100000;
		logarithm_table[2436] = 14'b0000100_0100000;
		logarithm_table[2437] = 14'b0000100_0100000;
		logarithm_table[2438] = 14'b0000100_0100000;
		logarithm_table[2439] = 14'b0000100_0100000;
		logarithm_table[2440] = 14'b0000100_0100000;
		logarithm_table[2441] = 14'b0000100_0100000;
		logarithm_table[2442] = 14'b0000100_0100000;
		logarithm_table[2443] = 14'b0000100_0100001;
		logarithm_table[2444] = 14'b0000100_0100001;
		logarithm_table[2445] = 14'b0000100_0100001;
		logarithm_table[2446] = 14'b0000100_0100001;
		logarithm_table[2447] = 14'b0000100_0100001;
		logarithm_table[2448] = 14'b0000100_0100001;
		logarithm_table[2449] = 14'b0000100_0100001;
		logarithm_table[2450] = 14'b0000100_0100001;
		logarithm_table[2451] = 14'b0000100_0100001;
		logarithm_table[2452] = 14'b0000100_0100001;
		logarithm_table[2453] = 14'b0000100_0100001;
		logarithm_table[2454] = 14'b0000100_0100001;
		logarithm_table[2455] = 14'b0000100_0100001;
		logarithm_table[2456] = 14'b0000100_0100010;
		logarithm_table[2457] = 14'b0000100_0100010;
		logarithm_table[2458] = 14'b0000100_0100010;
		logarithm_table[2459] = 14'b0000100_0100010;
		logarithm_table[2460] = 14'b0000100_0100010;
		logarithm_table[2461] = 14'b0000100_0100010;
		logarithm_table[2462] = 14'b0000100_0100010;
		logarithm_table[2463] = 14'b0000100_0100010;
		logarithm_table[2464] = 14'b0000100_0100010;
		logarithm_table[2465] = 14'b0000100_0100010;
		logarithm_table[2466] = 14'b0000100_0100010;
		logarithm_table[2467] = 14'b0000100_0100010;
		logarithm_table[2468] = 14'b0000100_0100010;
		logarithm_table[2469] = 14'b0000100_0100011;
		logarithm_table[2470] = 14'b0000100_0100011;
		logarithm_table[2471] = 14'b0000100_0100011;
		logarithm_table[2472] = 14'b0000100_0100011;
		logarithm_table[2473] = 14'b0000100_0100011;
		logarithm_table[2474] = 14'b0000100_0100011;
		logarithm_table[2475] = 14'b0000100_0100011;
		logarithm_table[2476] = 14'b0000100_0100011;
		logarithm_table[2477] = 14'b0000100_0100011;
		logarithm_table[2478] = 14'b0000100_0100011;
		logarithm_table[2479] = 14'b0000100_0100011;
		logarithm_table[2480] = 14'b0000100_0100011;
		logarithm_table[2481] = 14'b0000100_0100011;
		logarithm_table[2482] = 14'b0000100_0100011;
		logarithm_table[2483] = 14'b0000100_0100100;
		logarithm_table[2484] = 14'b0000100_0100100;
		logarithm_table[2485] = 14'b0000100_0100100;
		logarithm_table[2486] = 14'b0000100_0100100;
		logarithm_table[2487] = 14'b0000100_0100100;
		logarithm_table[2488] = 14'b0000100_0100100;
		logarithm_table[2489] = 14'b0000100_0100100;
		logarithm_table[2490] = 14'b0000100_0100100;
		logarithm_table[2491] = 14'b0000100_0100100;
		logarithm_table[2492] = 14'b0000100_0100100;
		logarithm_table[2493] = 14'b0000100_0100100;
		logarithm_table[2494] = 14'b0000100_0100100;
		logarithm_table[2495] = 14'b0000100_0100100;
		logarithm_table[2496] = 14'b0000100_0100101;
		logarithm_table[2497] = 14'b0000100_0100101;
		logarithm_table[2498] = 14'b0000100_0100101;
		logarithm_table[2499] = 14'b0000100_0100101;
		logarithm_table[2500] = 14'b0000100_0100101;
		logarithm_table[2501] = 14'b0000100_0100101;
		logarithm_table[2502] = 14'b0000100_0100101;
		logarithm_table[2503] = 14'b0000100_0100101;
		logarithm_table[2504] = 14'b0000100_0100101;
		logarithm_table[2505] = 14'b0000100_0100101;
		logarithm_table[2506] = 14'b0000100_0100101;
		logarithm_table[2507] = 14'b0000100_0100101;
		logarithm_table[2508] = 14'b0000100_0100101;
		logarithm_table[2509] = 14'b0000100_0100101;
		logarithm_table[2510] = 14'b0000100_0100110;
		logarithm_table[2511] = 14'b0000100_0100110;
		logarithm_table[2512] = 14'b0000100_0100110;
		logarithm_table[2513] = 14'b0000100_0100110;
		logarithm_table[2514] = 14'b0000100_0100110;
		logarithm_table[2515] = 14'b0000100_0100110;
		logarithm_table[2516] = 14'b0000100_0100110;
		logarithm_table[2517] = 14'b0000100_0100110;
		logarithm_table[2518] = 14'b0000100_0100110;
		logarithm_table[2519] = 14'b0000100_0100110;
		logarithm_table[2520] = 14'b0000100_0100110;
		logarithm_table[2521] = 14'b0000100_0100110;
		logarithm_table[2522] = 14'b0000100_0100110;
		logarithm_table[2523] = 14'b0000100_0100111;
		logarithm_table[2524] = 14'b0000100_0100111;
		logarithm_table[2525] = 14'b0000100_0100111;
		logarithm_table[2526] = 14'b0000100_0100111;
		logarithm_table[2527] = 14'b0000100_0100111;
		logarithm_table[2528] = 14'b0000100_0100111;
		logarithm_table[2529] = 14'b0000100_0100111;
		logarithm_table[2530] = 14'b0000100_0100111;
		logarithm_table[2531] = 14'b0000100_0100111;
		logarithm_table[2532] = 14'b0000100_0100111;
		logarithm_table[2533] = 14'b0000100_0100111;
		logarithm_table[2534] = 14'b0000100_0100111;
		logarithm_table[2535] = 14'b0000100_0100111;
		logarithm_table[2536] = 14'b0000100_0100111;
		logarithm_table[2537] = 14'b0000100_0101000;
		logarithm_table[2538] = 14'b0000100_0101000;
		logarithm_table[2539] = 14'b0000100_0101000;
		logarithm_table[2540] = 14'b0000100_0101000;
		logarithm_table[2541] = 14'b0000100_0101000;
		logarithm_table[2542] = 14'b0000100_0101000;
		logarithm_table[2543] = 14'b0000100_0101000;
		logarithm_table[2544] = 14'b0000100_0101000;
		logarithm_table[2545] = 14'b0000100_0101000;
		logarithm_table[2546] = 14'b0000100_0101000;
		logarithm_table[2547] = 14'b0000100_0101000;
		logarithm_table[2548] = 14'b0000100_0101000;
		logarithm_table[2549] = 14'b0000100_0101000;
		logarithm_table[2550] = 14'b0000100_0101000;
		logarithm_table[2551] = 14'b0000100_0101001;
		logarithm_table[2552] = 14'b0000100_0101001;
		logarithm_table[2553] = 14'b0000100_0101001;
		logarithm_table[2554] = 14'b0000100_0101001;
		logarithm_table[2555] = 14'b0000100_0101001;
		logarithm_table[2556] = 14'b0000100_0101001;
		logarithm_table[2557] = 14'b0000100_0101001;
		logarithm_table[2558] = 14'b0000100_0101001;
		logarithm_table[2559] = 14'b0000100_0101001;
		logarithm_table[2560] = 14'b0000100_0101001;
		logarithm_table[2561] = 14'b0000100_0101001;
		logarithm_table[2562] = 14'b0000100_0101001;
		logarithm_table[2563] = 14'b0000100_0101001;
		logarithm_table[2564] = 14'b0000100_0101001;
		logarithm_table[2565] = 14'b0000100_0101010;
		logarithm_table[2566] = 14'b0000100_0101010;
		logarithm_table[2567] = 14'b0000100_0101010;
		logarithm_table[2568] = 14'b0000100_0101010;
		logarithm_table[2569] = 14'b0000100_0101010;
		logarithm_table[2570] = 14'b0000100_0101010;
		logarithm_table[2571] = 14'b0000100_0101010;
		logarithm_table[2572] = 14'b0000100_0101010;
		logarithm_table[2573] = 14'b0000100_0101010;
		logarithm_table[2574] = 14'b0000100_0101010;
		logarithm_table[2575] = 14'b0000100_0101010;
		logarithm_table[2576] = 14'b0000100_0101010;
		logarithm_table[2577] = 14'b0000100_0101010;
		logarithm_table[2578] = 14'b0000100_0101011;
		logarithm_table[2579] = 14'b0000100_0101011;
		logarithm_table[2580] = 14'b0000100_0101011;
		logarithm_table[2581] = 14'b0000100_0101011;
		logarithm_table[2582] = 14'b0000100_0101011;
		logarithm_table[2583] = 14'b0000100_0101011;
		logarithm_table[2584] = 14'b0000100_0101011;
		logarithm_table[2585] = 14'b0000100_0101011;
		logarithm_table[2586] = 14'b0000100_0101011;
		logarithm_table[2587] = 14'b0000100_0101011;
		logarithm_table[2588] = 14'b0000100_0101011;
		logarithm_table[2589] = 14'b0000100_0101011;
		logarithm_table[2590] = 14'b0000100_0101011;
		logarithm_table[2591] = 14'b0000100_0101011;
		logarithm_table[2592] = 14'b0000100_0101100;
		logarithm_table[2593] = 14'b0000100_0101100;
		logarithm_table[2594] = 14'b0000100_0101100;
		logarithm_table[2595] = 14'b0000100_0101100;
		logarithm_table[2596] = 14'b0000100_0101100;
		logarithm_table[2597] = 14'b0000100_0101100;
		logarithm_table[2598] = 14'b0000100_0101100;
		logarithm_table[2599] = 14'b0000100_0101100;
		logarithm_table[2600] = 14'b0000100_0101100;
		logarithm_table[2601] = 14'b0000100_0101100;
		logarithm_table[2602] = 14'b0000100_0101100;
		logarithm_table[2603] = 14'b0000100_0101100;
		logarithm_table[2604] = 14'b0000100_0101100;
		logarithm_table[2605] = 14'b0000100_0101100;
		logarithm_table[2606] = 14'b0000100_0101100;
		logarithm_table[2607] = 14'b0000100_0101101;
		logarithm_table[2608] = 14'b0000100_0101101;
		logarithm_table[2609] = 14'b0000100_0101101;
		logarithm_table[2610] = 14'b0000100_0101101;
		logarithm_table[2611] = 14'b0000100_0101101;
		logarithm_table[2612] = 14'b0000100_0101101;
		logarithm_table[2613] = 14'b0000100_0101101;
		logarithm_table[2614] = 14'b0000100_0101101;
		logarithm_table[2615] = 14'b0000100_0101101;
		logarithm_table[2616] = 14'b0000100_0101101;
		logarithm_table[2617] = 14'b0000100_0101101;
		logarithm_table[2618] = 14'b0000100_0101101;
		logarithm_table[2619] = 14'b0000100_0101101;
		logarithm_table[2620] = 14'b0000100_0101101;
		logarithm_table[2621] = 14'b0000100_0101110;
		logarithm_table[2622] = 14'b0000100_0101110;
		logarithm_table[2623] = 14'b0000100_0101110;
		logarithm_table[2624] = 14'b0000100_0101110;
		logarithm_table[2625] = 14'b0000100_0101110;
		logarithm_table[2626] = 14'b0000100_0101110;
		logarithm_table[2627] = 14'b0000100_0101110;
		logarithm_table[2628] = 14'b0000100_0101110;
		logarithm_table[2629] = 14'b0000100_0101110;
		logarithm_table[2630] = 14'b0000100_0101110;
		logarithm_table[2631] = 14'b0000100_0101110;
		logarithm_table[2632] = 14'b0000100_0101110;
		logarithm_table[2633] = 14'b0000100_0101110;
		logarithm_table[2634] = 14'b0000100_0101110;
		logarithm_table[2635] = 14'b0000100_0101111;
		logarithm_table[2636] = 14'b0000100_0101111;
		logarithm_table[2637] = 14'b0000100_0101111;
		logarithm_table[2638] = 14'b0000100_0101111;
		logarithm_table[2639] = 14'b0000100_0101111;
		logarithm_table[2640] = 14'b0000100_0101111;
		logarithm_table[2641] = 14'b0000100_0101111;
		logarithm_table[2642] = 14'b0000100_0101111;
		logarithm_table[2643] = 14'b0000100_0101111;
		logarithm_table[2644] = 14'b0000100_0101111;
		logarithm_table[2645] = 14'b0000100_0101111;
		logarithm_table[2646] = 14'b0000100_0101111;
		logarithm_table[2647] = 14'b0000100_0101111;
		logarithm_table[2648] = 14'b0000100_0101111;
		logarithm_table[2649] = 14'b0000100_0110000;
		logarithm_table[2650] = 14'b0000100_0110000;
		logarithm_table[2651] = 14'b0000100_0110000;
		logarithm_table[2652] = 14'b0000100_0110000;
		logarithm_table[2653] = 14'b0000100_0110000;
		logarithm_table[2654] = 14'b0000100_0110000;
		logarithm_table[2655] = 14'b0000100_0110000;
		logarithm_table[2656] = 14'b0000100_0110000;
		logarithm_table[2657] = 14'b0000100_0110000;
		logarithm_table[2658] = 14'b0000100_0110000;
		logarithm_table[2659] = 14'b0000100_0110000;
		logarithm_table[2660] = 14'b0000100_0110000;
		logarithm_table[2661] = 14'b0000100_0110000;
		logarithm_table[2662] = 14'b0000100_0110000;
		logarithm_table[2663] = 14'b0000100_0110000;
		logarithm_table[2664] = 14'b0000100_0110001;
		logarithm_table[2665] = 14'b0000100_0110001;
		logarithm_table[2666] = 14'b0000100_0110001;
		logarithm_table[2667] = 14'b0000100_0110001;
		logarithm_table[2668] = 14'b0000100_0110001;
		logarithm_table[2669] = 14'b0000100_0110001;
		logarithm_table[2670] = 14'b0000100_0110001;
		logarithm_table[2671] = 14'b0000100_0110001;
		logarithm_table[2672] = 14'b0000100_0110001;
		logarithm_table[2673] = 14'b0000100_0110001;
		logarithm_table[2674] = 14'b0000100_0110001;
		logarithm_table[2675] = 14'b0000100_0110001;
		logarithm_table[2676] = 14'b0000100_0110001;
		logarithm_table[2677] = 14'b0000100_0110001;
		logarithm_table[2678] = 14'b0000100_0110010;
		logarithm_table[2679] = 14'b0000100_0110010;
		logarithm_table[2680] = 14'b0000100_0110010;
		logarithm_table[2681] = 14'b0000100_0110010;
		logarithm_table[2682] = 14'b0000100_0110010;
		logarithm_table[2683] = 14'b0000100_0110010;
		logarithm_table[2684] = 14'b0000100_0110010;
		logarithm_table[2685] = 14'b0000100_0110010;
		logarithm_table[2686] = 14'b0000100_0110010;
		logarithm_table[2687] = 14'b0000100_0110010;
		logarithm_table[2688] = 14'b0000100_0110010;
		logarithm_table[2689] = 14'b0000100_0110010;
		logarithm_table[2690] = 14'b0000100_0110010;
		logarithm_table[2691] = 14'b0000100_0110010;
		logarithm_table[2692] = 14'b0000100_0110010;
		logarithm_table[2693] = 14'b0000100_0110011;
		logarithm_table[2694] = 14'b0000100_0110011;
		logarithm_table[2695] = 14'b0000100_0110011;
		logarithm_table[2696] = 14'b0000100_0110011;
		logarithm_table[2697] = 14'b0000100_0110011;
		logarithm_table[2698] = 14'b0000100_0110011;
		logarithm_table[2699] = 14'b0000100_0110011;
		logarithm_table[2700] = 14'b0000100_0110011;
		logarithm_table[2701] = 14'b0000100_0110011;
		logarithm_table[2702] = 14'b0000100_0110011;
		logarithm_table[2703] = 14'b0000100_0110011;
		logarithm_table[2704] = 14'b0000100_0110011;
		logarithm_table[2705] = 14'b0000100_0110011;
		logarithm_table[2706] = 14'b0000100_0110011;
		logarithm_table[2707] = 14'b0000100_0110100;
		logarithm_table[2708] = 14'b0000100_0110100;
		logarithm_table[2709] = 14'b0000100_0110100;
		logarithm_table[2710] = 14'b0000100_0110100;
		logarithm_table[2711] = 14'b0000100_0110100;
		logarithm_table[2712] = 14'b0000100_0110100;
		logarithm_table[2713] = 14'b0000100_0110100;
		logarithm_table[2714] = 14'b0000100_0110100;
		logarithm_table[2715] = 14'b0000100_0110100;
		logarithm_table[2716] = 14'b0000100_0110100;
		logarithm_table[2717] = 14'b0000100_0110100;
		logarithm_table[2718] = 14'b0000100_0110100;
		logarithm_table[2719] = 14'b0000100_0110100;
		logarithm_table[2720] = 14'b0000100_0110100;
		logarithm_table[2721] = 14'b0000100_0110100;
		logarithm_table[2722] = 14'b0000100_0110101;
		logarithm_table[2723] = 14'b0000100_0110101;
		logarithm_table[2724] = 14'b0000100_0110101;
		logarithm_table[2725] = 14'b0000100_0110101;
		logarithm_table[2726] = 14'b0000100_0110101;
		logarithm_table[2727] = 14'b0000100_0110101;
		logarithm_table[2728] = 14'b0000100_0110101;
		logarithm_table[2729] = 14'b0000100_0110101;
		logarithm_table[2730] = 14'b0000100_0110101;
		logarithm_table[2731] = 14'b0000100_0110101;
		logarithm_table[2732] = 14'b0000100_0110101;
		logarithm_table[2733] = 14'b0000100_0110101;
		logarithm_table[2734] = 14'b0000100_0110101;
		logarithm_table[2735] = 14'b0000100_0110101;
		logarithm_table[2736] = 14'b0000100_0110101;
		logarithm_table[2737] = 14'b0000100_0110110;
		logarithm_table[2738] = 14'b0000100_0110110;
		logarithm_table[2739] = 14'b0000100_0110110;
		logarithm_table[2740] = 14'b0000100_0110110;
		logarithm_table[2741] = 14'b0000100_0110110;
		logarithm_table[2742] = 14'b0000100_0110110;
		logarithm_table[2743] = 14'b0000100_0110110;
		logarithm_table[2744] = 14'b0000100_0110110;
		logarithm_table[2745] = 14'b0000100_0110110;
		logarithm_table[2746] = 14'b0000100_0110110;
		logarithm_table[2747] = 14'b0000100_0110110;
		logarithm_table[2748] = 14'b0000100_0110110;
		logarithm_table[2749] = 14'b0000100_0110110;
		logarithm_table[2750] = 14'b0000100_0110110;
		logarithm_table[2751] = 14'b0000100_0110110;
		logarithm_table[2752] = 14'b0000100_0110111;
		logarithm_table[2753] = 14'b0000100_0110111;
		logarithm_table[2754] = 14'b0000100_0110111;
		logarithm_table[2755] = 14'b0000100_0110111;
		logarithm_table[2756] = 14'b0000100_0110111;
		logarithm_table[2757] = 14'b0000100_0110111;
		logarithm_table[2758] = 14'b0000100_0110111;
		logarithm_table[2759] = 14'b0000100_0110111;
		logarithm_table[2760] = 14'b0000100_0110111;
		logarithm_table[2761] = 14'b0000100_0110111;
		logarithm_table[2762] = 14'b0000100_0110111;
		logarithm_table[2763] = 14'b0000100_0110111;
		logarithm_table[2764] = 14'b0000100_0110111;
		logarithm_table[2765] = 14'b0000100_0110111;
		logarithm_table[2766] = 14'b0000100_0110111;
		logarithm_table[2767] = 14'b0000100_0111000;
		logarithm_table[2768] = 14'b0000100_0111000;
		logarithm_table[2769] = 14'b0000100_0111000;
		logarithm_table[2770] = 14'b0000100_0111000;
		logarithm_table[2771] = 14'b0000100_0111000;
		logarithm_table[2772] = 14'b0000100_0111000;
		logarithm_table[2773] = 14'b0000100_0111000;
		logarithm_table[2774] = 14'b0000100_0111000;
		logarithm_table[2775] = 14'b0000100_0111000;
		logarithm_table[2776] = 14'b0000100_0111000;
		logarithm_table[2777] = 14'b0000100_0111000;
		logarithm_table[2778] = 14'b0000100_0111000;
		logarithm_table[2779] = 14'b0000100_0111000;
		logarithm_table[2780] = 14'b0000100_0111000;
		logarithm_table[2781] = 14'b0000100_0111000;
		logarithm_table[2782] = 14'b0000100_0111001;
		logarithm_table[2783] = 14'b0000100_0111001;
		logarithm_table[2784] = 14'b0000100_0111001;
		logarithm_table[2785] = 14'b0000100_0111001;
		logarithm_table[2786] = 14'b0000100_0111001;
		logarithm_table[2787] = 14'b0000100_0111001;
		logarithm_table[2788] = 14'b0000100_0111001;
		logarithm_table[2789] = 14'b0000100_0111001;
		logarithm_table[2790] = 14'b0000100_0111001;
		logarithm_table[2791] = 14'b0000100_0111001;
		logarithm_table[2792] = 14'b0000100_0111001;
		logarithm_table[2793] = 14'b0000100_0111001;
		logarithm_table[2794] = 14'b0000100_0111001;
		logarithm_table[2795] = 14'b0000100_0111001;
		logarithm_table[2796] = 14'b0000100_0111001;
		logarithm_table[2797] = 14'b0000100_0111010;
		logarithm_table[2798] = 14'b0000100_0111010;
		logarithm_table[2799] = 14'b0000100_0111010;
		logarithm_table[2800] = 14'b0000100_0111010;
		logarithm_table[2801] = 14'b0000100_0111010;
		logarithm_table[2802] = 14'b0000100_0111010;
		logarithm_table[2803] = 14'b0000100_0111010;
		logarithm_table[2804] = 14'b0000100_0111010;
		logarithm_table[2805] = 14'b0000100_0111010;
		logarithm_table[2806] = 14'b0000100_0111010;
		logarithm_table[2807] = 14'b0000100_0111010;
		logarithm_table[2808] = 14'b0000100_0111010;
		logarithm_table[2809] = 14'b0000100_0111010;
		logarithm_table[2810] = 14'b0000100_0111010;
		logarithm_table[2811] = 14'b0000100_0111010;
		logarithm_table[2812] = 14'b0000100_0111011;
		logarithm_table[2813] = 14'b0000100_0111011;
		logarithm_table[2814] = 14'b0000100_0111011;
		logarithm_table[2815] = 14'b0000100_0111011;
		logarithm_table[2816] = 14'b0000100_0111011;
		logarithm_table[2817] = 14'b0000100_0111011;
		logarithm_table[2818] = 14'b0000100_0111011;
		logarithm_table[2819] = 14'b0000100_0111011;
		logarithm_table[2820] = 14'b0000100_0111011;
		logarithm_table[2821] = 14'b0000100_0111011;
		logarithm_table[2822] = 14'b0000100_0111011;
		logarithm_table[2823] = 14'b0000100_0111011;
		logarithm_table[2824] = 14'b0000100_0111011;
		logarithm_table[2825] = 14'b0000100_0111011;
		logarithm_table[2826] = 14'b0000100_0111011;
		logarithm_table[2827] = 14'b0000100_0111100;
		logarithm_table[2828] = 14'b0000100_0111100;
		logarithm_table[2829] = 14'b0000100_0111100;
		logarithm_table[2830] = 14'b0000100_0111100;
		logarithm_table[2831] = 14'b0000100_0111100;
		logarithm_table[2832] = 14'b0000100_0111100;
		logarithm_table[2833] = 14'b0000100_0111100;
		logarithm_table[2834] = 14'b0000100_0111100;
		logarithm_table[2835] = 14'b0000100_0111100;
		logarithm_table[2836] = 14'b0000100_0111100;
		logarithm_table[2837] = 14'b0000100_0111100;
		logarithm_table[2838] = 14'b0000100_0111100;
		logarithm_table[2839] = 14'b0000100_0111100;
		logarithm_table[2840] = 14'b0000100_0111100;
		logarithm_table[2841] = 14'b0000100_0111100;
		logarithm_table[2842] = 14'b0000100_0111101;
		logarithm_table[2843] = 14'b0000100_0111101;
		logarithm_table[2844] = 14'b0000100_0111101;
		logarithm_table[2845] = 14'b0000100_0111101;
		logarithm_table[2846] = 14'b0000100_0111101;
		logarithm_table[2847] = 14'b0000100_0111101;
		logarithm_table[2848] = 14'b0000100_0111101;
		logarithm_table[2849] = 14'b0000100_0111101;
		logarithm_table[2850] = 14'b0000100_0111101;
		logarithm_table[2851] = 14'b0000100_0111101;
		logarithm_table[2852] = 14'b0000100_0111101;
		logarithm_table[2853] = 14'b0000100_0111101;
		logarithm_table[2854] = 14'b0000100_0111101;
		logarithm_table[2855] = 14'b0000100_0111101;
		logarithm_table[2856] = 14'b0000100_0111101;
		logarithm_table[2857] = 14'b0000100_0111101;
		logarithm_table[2858] = 14'b0000100_0111110;
		logarithm_table[2859] = 14'b0000100_0111110;
		logarithm_table[2860] = 14'b0000100_0111110;
		logarithm_table[2861] = 14'b0000100_0111110;
		logarithm_table[2862] = 14'b0000100_0111110;
		logarithm_table[2863] = 14'b0000100_0111110;
		logarithm_table[2864] = 14'b0000100_0111110;
		logarithm_table[2865] = 14'b0000100_0111110;
		logarithm_table[2866] = 14'b0000100_0111110;
		logarithm_table[2867] = 14'b0000100_0111110;
		logarithm_table[2868] = 14'b0000100_0111110;
		logarithm_table[2869] = 14'b0000100_0111110;
		logarithm_table[2870] = 14'b0000100_0111110;
		logarithm_table[2871] = 14'b0000100_0111110;
		logarithm_table[2872] = 14'b0000100_0111110;
		logarithm_table[2873] = 14'b0000100_0111111;
		logarithm_table[2874] = 14'b0000100_0111111;
		logarithm_table[2875] = 14'b0000100_0111111;
		logarithm_table[2876] = 14'b0000100_0111111;
		logarithm_table[2877] = 14'b0000100_0111111;
		logarithm_table[2878] = 14'b0000100_0111111;
		logarithm_table[2879] = 14'b0000100_0111111;
		logarithm_table[2880] = 14'b0000100_0111111;
		logarithm_table[2881] = 14'b0000100_0111111;
		logarithm_table[2882] = 14'b0000100_0111111;
		logarithm_table[2883] = 14'b0000100_0111111;
		logarithm_table[2884] = 14'b0000100_0111111;
		logarithm_table[2885] = 14'b0000100_0111111;
		logarithm_table[2886] = 14'b0000100_0111111;
		logarithm_table[2887] = 14'b0000100_0111111;
		logarithm_table[2888] = 14'b0000100_0111111;
		logarithm_table[2889] = 14'b0000100_1000000;
		logarithm_table[2890] = 14'b0000100_1000000;
		logarithm_table[2891] = 14'b0000100_1000000;
		logarithm_table[2892] = 14'b0000100_1000000;
		logarithm_table[2893] = 14'b0000100_1000000;
		logarithm_table[2894] = 14'b0000100_1000000;
		logarithm_table[2895] = 14'b0000100_1000000;
		logarithm_table[2896] = 14'b0000100_1000000;
		logarithm_table[2897] = 14'b0000100_1000000;
		logarithm_table[2898] = 14'b0000100_1000000;
		logarithm_table[2899] = 14'b0000100_1000000;
		logarithm_table[2900] = 14'b0000100_1000000;
		logarithm_table[2901] = 14'b0000100_1000000;
		logarithm_table[2902] = 14'b0000100_1000000;
		logarithm_table[2903] = 14'b0000100_1000000;
		logarithm_table[2904] = 14'b0000100_1000000;
		logarithm_table[2905] = 14'b0000100_1000001;
		logarithm_table[2906] = 14'b0000100_1000001;
		logarithm_table[2907] = 14'b0000100_1000001;
		logarithm_table[2908] = 14'b0000100_1000001;
		logarithm_table[2909] = 14'b0000100_1000001;
		logarithm_table[2910] = 14'b0000100_1000001;
		logarithm_table[2911] = 14'b0000100_1000001;
		logarithm_table[2912] = 14'b0000100_1000001;
		logarithm_table[2913] = 14'b0000100_1000001;
		logarithm_table[2914] = 14'b0000100_1000001;
		logarithm_table[2915] = 14'b0000100_1000001;
		logarithm_table[2916] = 14'b0000100_1000001;
		logarithm_table[2917] = 14'b0000100_1000001;
		logarithm_table[2918] = 14'b0000100_1000001;
		logarithm_table[2919] = 14'b0000100_1000001;
		logarithm_table[2920] = 14'b0000100_1000010;
		logarithm_table[2921] = 14'b0000100_1000010;
		logarithm_table[2922] = 14'b0000100_1000010;
		logarithm_table[2923] = 14'b0000100_1000010;
		logarithm_table[2924] = 14'b0000100_1000010;
		logarithm_table[2925] = 14'b0000100_1000010;
		logarithm_table[2926] = 14'b0000100_1000010;
		logarithm_table[2927] = 14'b0000100_1000010;
		logarithm_table[2928] = 14'b0000100_1000010;
		logarithm_table[2929] = 14'b0000100_1000010;
		logarithm_table[2930] = 14'b0000100_1000010;
		logarithm_table[2931] = 14'b0000100_1000010;
		logarithm_table[2932] = 14'b0000100_1000010;
		logarithm_table[2933] = 14'b0000100_1000010;
		logarithm_table[2934] = 14'b0000100_1000010;
		logarithm_table[2935] = 14'b0000100_1000010;
		logarithm_table[2936] = 14'b0000100_1000011;
		logarithm_table[2937] = 14'b0000100_1000011;
		logarithm_table[2938] = 14'b0000100_1000011;
		logarithm_table[2939] = 14'b0000100_1000011;
		logarithm_table[2940] = 14'b0000100_1000011;
		logarithm_table[2941] = 14'b0000100_1000011;
		logarithm_table[2942] = 14'b0000100_1000011;
		logarithm_table[2943] = 14'b0000100_1000011;
		logarithm_table[2944] = 14'b0000100_1000011;
		logarithm_table[2945] = 14'b0000100_1000011;
		logarithm_table[2946] = 14'b0000100_1000011;
		logarithm_table[2947] = 14'b0000100_1000011;
		logarithm_table[2948] = 14'b0000100_1000011;
		logarithm_table[2949] = 14'b0000100_1000011;
		logarithm_table[2950] = 14'b0000100_1000011;
		logarithm_table[2951] = 14'b0000100_1000011;
		logarithm_table[2952] = 14'b0000100_1000100;
		logarithm_table[2953] = 14'b0000100_1000100;
		logarithm_table[2954] = 14'b0000100_1000100;
		logarithm_table[2955] = 14'b0000100_1000100;
		logarithm_table[2956] = 14'b0000100_1000100;
		logarithm_table[2957] = 14'b0000100_1000100;
		logarithm_table[2958] = 14'b0000100_1000100;
		logarithm_table[2959] = 14'b0000100_1000100;
		logarithm_table[2960] = 14'b0000100_1000100;
		logarithm_table[2961] = 14'b0000100_1000100;
		logarithm_table[2962] = 14'b0000100_1000100;
		logarithm_table[2963] = 14'b0000100_1000100;
		logarithm_table[2964] = 14'b0000100_1000100;
		logarithm_table[2965] = 14'b0000100_1000100;
		logarithm_table[2966] = 14'b0000100_1000100;
		logarithm_table[2967] = 14'b0000100_1000100;
		logarithm_table[2968] = 14'b0000100_1000101;
		logarithm_table[2969] = 14'b0000100_1000101;
		logarithm_table[2970] = 14'b0000100_1000101;
		logarithm_table[2971] = 14'b0000100_1000101;
		logarithm_table[2972] = 14'b0000100_1000101;
		logarithm_table[2973] = 14'b0000100_1000101;
		logarithm_table[2974] = 14'b0000100_1000101;
		logarithm_table[2975] = 14'b0000100_1000101;
		logarithm_table[2976] = 14'b0000100_1000101;
		logarithm_table[2977] = 14'b0000100_1000101;
		logarithm_table[2978] = 14'b0000100_1000101;
		logarithm_table[2979] = 14'b0000100_1000101;
		logarithm_table[2980] = 14'b0000100_1000101;
		logarithm_table[2981] = 14'b0000100_1000101;
		logarithm_table[2982] = 14'b0000100_1000101;
		logarithm_table[2983] = 14'b0000100_1000101;
		logarithm_table[2984] = 14'b0000100_1000110;
		logarithm_table[2985] = 14'b0000100_1000110;
		logarithm_table[2986] = 14'b0000100_1000110;
		logarithm_table[2987] = 14'b0000100_1000110;
		logarithm_table[2988] = 14'b0000100_1000110;
		logarithm_table[2989] = 14'b0000100_1000110;
		logarithm_table[2990] = 14'b0000100_1000110;
		logarithm_table[2991] = 14'b0000100_1000110;
		logarithm_table[2992] = 14'b0000100_1000110;
		logarithm_table[2993] = 14'b0000100_1000110;
		logarithm_table[2994] = 14'b0000100_1000110;
		logarithm_table[2995] = 14'b0000100_1000110;
		logarithm_table[2996] = 14'b0000100_1000110;
		logarithm_table[2997] = 14'b0000100_1000110;
		logarithm_table[2998] = 14'b0000100_1000110;
		logarithm_table[2999] = 14'b0000100_1000110;
		logarithm_table[3000] = 14'b0000100_1000110;
		logarithm_table[3001] = 14'b0000100_1000111;
		logarithm_table[3002] = 14'b0000100_1000111;
		logarithm_table[3003] = 14'b0000100_1000111;
		logarithm_table[3004] = 14'b0000100_1000111;
		logarithm_table[3005] = 14'b0000100_1000111;
		logarithm_table[3006] = 14'b0000100_1000111;
		logarithm_table[3007] = 14'b0000100_1000111;
		logarithm_table[3008] = 14'b0000100_1000111;
		logarithm_table[3009] = 14'b0000100_1000111;
		logarithm_table[3010] = 14'b0000100_1000111;
		logarithm_table[3011] = 14'b0000100_1000111;
		logarithm_table[3012] = 14'b0000100_1000111;
		logarithm_table[3013] = 14'b0000100_1000111;
		logarithm_table[3014] = 14'b0000100_1000111;
		logarithm_table[3015] = 14'b0000100_1000111;
		logarithm_table[3016] = 14'b0000100_1000111;
		logarithm_table[3017] = 14'b0000100_1001000;
		logarithm_table[3018] = 14'b0000100_1001000;
		logarithm_table[3019] = 14'b0000100_1001000;
		logarithm_table[3020] = 14'b0000100_1001000;
		logarithm_table[3021] = 14'b0000100_1001000;
		logarithm_table[3022] = 14'b0000100_1001000;
		logarithm_table[3023] = 14'b0000100_1001000;
		logarithm_table[3024] = 14'b0000100_1001000;
		logarithm_table[3025] = 14'b0000100_1001000;
		logarithm_table[3026] = 14'b0000100_1001000;
		logarithm_table[3027] = 14'b0000100_1001000;
		logarithm_table[3028] = 14'b0000100_1001000;
		logarithm_table[3029] = 14'b0000100_1001000;
		logarithm_table[3030] = 14'b0000100_1001000;
		logarithm_table[3031] = 14'b0000100_1001000;
		logarithm_table[3032] = 14'b0000100_1001000;
		logarithm_table[3033] = 14'b0000100_1001001;
		logarithm_table[3034] = 14'b0000100_1001001;
		logarithm_table[3035] = 14'b0000100_1001001;
		logarithm_table[3036] = 14'b0000100_1001001;
		logarithm_table[3037] = 14'b0000100_1001001;
		logarithm_table[3038] = 14'b0000100_1001001;
		logarithm_table[3039] = 14'b0000100_1001001;
		logarithm_table[3040] = 14'b0000100_1001001;
		logarithm_table[3041] = 14'b0000100_1001001;
		logarithm_table[3042] = 14'b0000100_1001001;
		logarithm_table[3043] = 14'b0000100_1001001;
		logarithm_table[3044] = 14'b0000100_1001001;
		logarithm_table[3045] = 14'b0000100_1001001;
		logarithm_table[3046] = 14'b0000100_1001001;
		logarithm_table[3047] = 14'b0000100_1001001;
		logarithm_table[3048] = 14'b0000100_1001001;
		logarithm_table[3049] = 14'b0000100_1001001;
		logarithm_table[3050] = 14'b0000100_1001010;
		logarithm_table[3051] = 14'b0000100_1001010;
		logarithm_table[3052] = 14'b0000100_1001010;
		logarithm_table[3053] = 14'b0000100_1001010;
		logarithm_table[3054] = 14'b0000100_1001010;
		logarithm_table[3055] = 14'b0000100_1001010;
		logarithm_table[3056] = 14'b0000100_1001010;
		logarithm_table[3057] = 14'b0000100_1001010;
		logarithm_table[3058] = 14'b0000100_1001010;
		logarithm_table[3059] = 14'b0000100_1001010;
		logarithm_table[3060] = 14'b0000100_1001010;
		logarithm_table[3061] = 14'b0000100_1001010;
		logarithm_table[3062] = 14'b0000100_1001010;
		logarithm_table[3063] = 14'b0000100_1001010;
		logarithm_table[3064] = 14'b0000100_1001010;
		logarithm_table[3065] = 14'b0000100_1001010;
		logarithm_table[3066] = 14'b0000100_1001011;
		logarithm_table[3067] = 14'b0000100_1001011;
		logarithm_table[3068] = 14'b0000100_1001011;
		logarithm_table[3069] = 14'b0000100_1001011;
		logarithm_table[3070] = 14'b0000100_1001011;
		logarithm_table[3071] = 14'b0000100_1001011;
		logarithm_table[3072] = 14'b0000100_1001011;
		logarithm_table[3073] = 14'b0000100_1001011;
		logarithm_table[3074] = 14'b0000100_1001011;
		logarithm_table[3075] = 14'b0000100_1001011;
		logarithm_table[3076] = 14'b0000100_1001011;
		logarithm_table[3077] = 14'b0000100_1001011;
		logarithm_table[3078] = 14'b0000100_1001011;
		logarithm_table[3079] = 14'b0000100_1001011;
		logarithm_table[3080] = 14'b0000100_1001011;
		logarithm_table[3081] = 14'b0000100_1001011;
		logarithm_table[3082] = 14'b0000100_1001011;
		logarithm_table[3083] = 14'b0000100_1001100;
		logarithm_table[3084] = 14'b0000100_1001100;
		logarithm_table[3085] = 14'b0000100_1001100;
		logarithm_table[3086] = 14'b0000100_1001100;
		logarithm_table[3087] = 14'b0000100_1001100;
		logarithm_table[3088] = 14'b0000100_1001100;
		logarithm_table[3089] = 14'b0000100_1001100;
		logarithm_table[3090] = 14'b0000100_1001100;
		logarithm_table[3091] = 14'b0000100_1001100;
		logarithm_table[3092] = 14'b0000100_1001100;
		logarithm_table[3093] = 14'b0000100_1001100;
		logarithm_table[3094] = 14'b0000100_1001100;
		logarithm_table[3095] = 14'b0000100_1001100;
		logarithm_table[3096] = 14'b0000100_1001100;
		logarithm_table[3097] = 14'b0000100_1001100;
		logarithm_table[3098] = 14'b0000100_1001100;
		logarithm_table[3099] = 14'b0000100_1001100;
		logarithm_table[3100] = 14'b0000100_1001101;
		logarithm_table[3101] = 14'b0000100_1001101;
		logarithm_table[3102] = 14'b0000100_1001101;
		logarithm_table[3103] = 14'b0000100_1001101;
		logarithm_table[3104] = 14'b0000100_1001101;
		logarithm_table[3105] = 14'b0000100_1001101;
		logarithm_table[3106] = 14'b0000100_1001101;
		logarithm_table[3107] = 14'b0000100_1001101;
		logarithm_table[3108] = 14'b0000100_1001101;
		logarithm_table[3109] = 14'b0000100_1001101;
		logarithm_table[3110] = 14'b0000100_1001101;
		logarithm_table[3111] = 14'b0000100_1001101;
		logarithm_table[3112] = 14'b0000100_1001101;
		logarithm_table[3113] = 14'b0000100_1001101;
		logarithm_table[3114] = 14'b0000100_1001101;
		logarithm_table[3115] = 14'b0000100_1001101;
		logarithm_table[3116] = 14'b0000100_1001110;
		logarithm_table[3117] = 14'b0000100_1001110;
		logarithm_table[3118] = 14'b0000100_1001110;
		logarithm_table[3119] = 14'b0000100_1001110;
		logarithm_table[3120] = 14'b0000100_1001110;
		logarithm_table[3121] = 14'b0000100_1001110;
		logarithm_table[3122] = 14'b0000100_1001110;
		logarithm_table[3123] = 14'b0000100_1001110;
		logarithm_table[3124] = 14'b0000100_1001110;
		logarithm_table[3125] = 14'b0000100_1001110;
		logarithm_table[3126] = 14'b0000100_1001110;
		logarithm_table[3127] = 14'b0000100_1001110;
		logarithm_table[3128] = 14'b0000100_1001110;
		logarithm_table[3129] = 14'b0000100_1001110;
		logarithm_table[3130] = 14'b0000100_1001110;
		logarithm_table[3131] = 14'b0000100_1001110;
		logarithm_table[3132] = 14'b0000100_1001110;
		logarithm_table[3133] = 14'b0000100_1001111;
		logarithm_table[3134] = 14'b0000100_1001111;
		logarithm_table[3135] = 14'b0000100_1001111;
		logarithm_table[3136] = 14'b0000100_1001111;
		logarithm_table[3137] = 14'b0000100_1001111;
		logarithm_table[3138] = 14'b0000100_1001111;
		logarithm_table[3139] = 14'b0000100_1001111;
		logarithm_table[3140] = 14'b0000100_1001111;
		logarithm_table[3141] = 14'b0000100_1001111;
		logarithm_table[3142] = 14'b0000100_1001111;
		logarithm_table[3143] = 14'b0000100_1001111;
		logarithm_table[3144] = 14'b0000100_1001111;
		logarithm_table[3145] = 14'b0000100_1001111;
		logarithm_table[3146] = 14'b0000100_1001111;
		logarithm_table[3147] = 14'b0000100_1001111;
		logarithm_table[3148] = 14'b0000100_1001111;
		logarithm_table[3149] = 14'b0000100_1001111;
		logarithm_table[3150] = 14'b0000100_1010000;
		logarithm_table[3151] = 14'b0000100_1010000;
		logarithm_table[3152] = 14'b0000100_1010000;
		logarithm_table[3153] = 14'b0000100_1010000;
		logarithm_table[3154] = 14'b0000100_1010000;
		logarithm_table[3155] = 14'b0000100_1010000;
		logarithm_table[3156] = 14'b0000100_1010000;
		logarithm_table[3157] = 14'b0000100_1010000;
		logarithm_table[3158] = 14'b0000100_1010000;
		logarithm_table[3159] = 14'b0000100_1010000;
		logarithm_table[3160] = 14'b0000100_1010000;
		logarithm_table[3161] = 14'b0000100_1010000;
		logarithm_table[3162] = 14'b0000100_1010000;
		logarithm_table[3163] = 14'b0000100_1010000;
		logarithm_table[3164] = 14'b0000100_1010000;
		logarithm_table[3165] = 14'b0000100_1010000;
		logarithm_table[3166] = 14'b0000100_1010000;
		logarithm_table[3167] = 14'b0000100_1010000;
		logarithm_table[3168] = 14'b0000100_1010001;
		logarithm_table[3169] = 14'b0000100_1010001;
		logarithm_table[3170] = 14'b0000100_1010001;
		logarithm_table[3171] = 14'b0000100_1010001;
		logarithm_table[3172] = 14'b0000100_1010001;
		logarithm_table[3173] = 14'b0000100_1010001;
		logarithm_table[3174] = 14'b0000100_1010001;
		logarithm_table[3175] = 14'b0000100_1010001;
		logarithm_table[3176] = 14'b0000100_1010001;
		logarithm_table[3177] = 14'b0000100_1010001;
		logarithm_table[3178] = 14'b0000100_1010001;
		logarithm_table[3179] = 14'b0000100_1010001;
		logarithm_table[3180] = 14'b0000100_1010001;
		logarithm_table[3181] = 14'b0000100_1010001;
		logarithm_table[3182] = 14'b0000100_1010001;
		logarithm_table[3183] = 14'b0000100_1010001;
		logarithm_table[3184] = 14'b0000100_1010001;
		logarithm_table[3185] = 14'b0000100_1010010;
		logarithm_table[3186] = 14'b0000100_1010010;
		logarithm_table[3187] = 14'b0000100_1010010;
		logarithm_table[3188] = 14'b0000100_1010010;
		logarithm_table[3189] = 14'b0000100_1010010;
		logarithm_table[3190] = 14'b0000100_1010010;
		logarithm_table[3191] = 14'b0000100_1010010;
		logarithm_table[3192] = 14'b0000100_1010010;
		logarithm_table[3193] = 14'b0000100_1010010;
		logarithm_table[3194] = 14'b0000100_1010010;
		logarithm_table[3195] = 14'b0000100_1010010;
		logarithm_table[3196] = 14'b0000100_1010010;
		logarithm_table[3197] = 14'b0000100_1010010;
		logarithm_table[3198] = 14'b0000100_1010010;
		logarithm_table[3199] = 14'b0000100_1010010;
		logarithm_table[3200] = 14'b0000100_1010010;
		logarithm_table[3201] = 14'b0000100_1010010;
		logarithm_table[3202] = 14'b0000100_1010011;
		logarithm_table[3203] = 14'b0000100_1010011;
		logarithm_table[3204] = 14'b0000100_1010011;
		logarithm_table[3205] = 14'b0000100_1010011;
		logarithm_table[3206] = 14'b0000100_1010011;
		logarithm_table[3207] = 14'b0000100_1010011;
		logarithm_table[3208] = 14'b0000100_1010011;
		logarithm_table[3209] = 14'b0000100_1010011;
		logarithm_table[3210] = 14'b0000100_1010011;
		logarithm_table[3211] = 14'b0000100_1010011;
		logarithm_table[3212] = 14'b0000100_1010011;
		logarithm_table[3213] = 14'b0000100_1010011;
		logarithm_table[3214] = 14'b0000100_1010011;
		logarithm_table[3215] = 14'b0000100_1010011;
		logarithm_table[3216] = 14'b0000100_1010011;
		logarithm_table[3217] = 14'b0000100_1010011;
		logarithm_table[3218] = 14'b0000100_1010011;
		logarithm_table[3219] = 14'b0000100_1010100;
		logarithm_table[3220] = 14'b0000100_1010100;
		logarithm_table[3221] = 14'b0000100_1010100;
		logarithm_table[3222] = 14'b0000100_1010100;
		logarithm_table[3223] = 14'b0000100_1010100;
		logarithm_table[3224] = 14'b0000100_1010100;
		logarithm_table[3225] = 14'b0000100_1010100;
		logarithm_table[3226] = 14'b0000100_1010100;
		logarithm_table[3227] = 14'b0000100_1010100;
		logarithm_table[3228] = 14'b0000100_1010100;
		logarithm_table[3229] = 14'b0000100_1010100;
		logarithm_table[3230] = 14'b0000100_1010100;
		logarithm_table[3231] = 14'b0000100_1010100;
		logarithm_table[3232] = 14'b0000100_1010100;
		logarithm_table[3233] = 14'b0000100_1010100;
		logarithm_table[3234] = 14'b0000100_1010100;
		logarithm_table[3235] = 14'b0000100_1010100;
		logarithm_table[3236] = 14'b0000100_1010100;
		logarithm_table[3237] = 14'b0000100_1010101;
		logarithm_table[3238] = 14'b0000100_1010101;
		logarithm_table[3239] = 14'b0000100_1010101;
		logarithm_table[3240] = 14'b0000100_1010101;
		logarithm_table[3241] = 14'b0000100_1010101;
		logarithm_table[3242] = 14'b0000100_1010101;
		logarithm_table[3243] = 14'b0000100_1010101;
		logarithm_table[3244] = 14'b0000100_1010101;
		logarithm_table[3245] = 14'b0000100_1010101;
		logarithm_table[3246] = 14'b0000100_1010101;
		logarithm_table[3247] = 14'b0000100_1010101;
		logarithm_table[3248] = 14'b0000100_1010101;
		logarithm_table[3249] = 14'b0000100_1010101;
		logarithm_table[3250] = 14'b0000100_1010101;
		logarithm_table[3251] = 14'b0000100_1010101;
		logarithm_table[3252] = 14'b0000100_1010101;
		logarithm_table[3253] = 14'b0000100_1010101;
		logarithm_table[3254] = 14'b0000100_1010110;
		logarithm_table[3255] = 14'b0000100_1010110;
		logarithm_table[3256] = 14'b0000100_1010110;
		logarithm_table[3257] = 14'b0000100_1010110;
		logarithm_table[3258] = 14'b0000100_1010110;
		logarithm_table[3259] = 14'b0000100_1010110;
		logarithm_table[3260] = 14'b0000100_1010110;
		logarithm_table[3261] = 14'b0000100_1010110;
		logarithm_table[3262] = 14'b0000100_1010110;
		logarithm_table[3263] = 14'b0000100_1010110;
		logarithm_table[3264] = 14'b0000100_1010110;
		logarithm_table[3265] = 14'b0000100_1010110;
		logarithm_table[3266] = 14'b0000100_1010110;
		logarithm_table[3267] = 14'b0000100_1010110;
		logarithm_table[3268] = 14'b0000100_1010110;
		logarithm_table[3269] = 14'b0000100_1010110;
		logarithm_table[3270] = 14'b0000100_1010110;
		logarithm_table[3271] = 14'b0000100_1010110;
		logarithm_table[3272] = 14'b0000100_1010111;
		logarithm_table[3273] = 14'b0000100_1010111;
		logarithm_table[3274] = 14'b0000100_1010111;
		logarithm_table[3275] = 14'b0000100_1010111;
		logarithm_table[3276] = 14'b0000100_1010111;
		logarithm_table[3277] = 14'b0000100_1010111;
		logarithm_table[3278] = 14'b0000100_1010111;
		logarithm_table[3279] = 14'b0000100_1010111;
		logarithm_table[3280] = 14'b0000100_1010111;
		logarithm_table[3281] = 14'b0000100_1010111;
		logarithm_table[3282] = 14'b0000100_1010111;
		logarithm_table[3283] = 14'b0000100_1010111;
		logarithm_table[3284] = 14'b0000100_1010111;
		logarithm_table[3285] = 14'b0000100_1010111;
		logarithm_table[3286] = 14'b0000100_1010111;
		logarithm_table[3287] = 14'b0000100_1010111;
		logarithm_table[3288] = 14'b0000100_1010111;
		logarithm_table[3289] = 14'b0000100_1010111;
		logarithm_table[3290] = 14'b0000100_1011000;
		logarithm_table[3291] = 14'b0000100_1011000;
		logarithm_table[3292] = 14'b0000100_1011000;
		logarithm_table[3293] = 14'b0000100_1011000;
		logarithm_table[3294] = 14'b0000100_1011000;
		logarithm_table[3295] = 14'b0000100_1011000;
		logarithm_table[3296] = 14'b0000100_1011000;
		logarithm_table[3297] = 14'b0000100_1011000;
		logarithm_table[3298] = 14'b0000100_1011000;
		logarithm_table[3299] = 14'b0000100_1011000;
		logarithm_table[3300] = 14'b0000100_1011000;
		logarithm_table[3301] = 14'b0000100_1011000;
		logarithm_table[3302] = 14'b0000100_1011000;
		logarithm_table[3303] = 14'b0000100_1011000;
		logarithm_table[3304] = 14'b0000100_1011000;
		logarithm_table[3305] = 14'b0000100_1011000;
		logarithm_table[3306] = 14'b0000100_1011000;
		logarithm_table[3307] = 14'b0000100_1011000;
		logarithm_table[3308] = 14'b0000100_1011001;
		logarithm_table[3309] = 14'b0000100_1011001;
		logarithm_table[3310] = 14'b0000100_1011001;
		logarithm_table[3311] = 14'b0000100_1011001;
		logarithm_table[3312] = 14'b0000100_1011001;
		logarithm_table[3313] = 14'b0000100_1011001;
		logarithm_table[3314] = 14'b0000100_1011001;
		logarithm_table[3315] = 14'b0000100_1011001;
		logarithm_table[3316] = 14'b0000100_1011001;
		logarithm_table[3317] = 14'b0000100_1011001;
		logarithm_table[3318] = 14'b0000100_1011001;
		logarithm_table[3319] = 14'b0000100_1011001;
		logarithm_table[3320] = 14'b0000100_1011001;
		logarithm_table[3321] = 14'b0000100_1011001;
		logarithm_table[3322] = 14'b0000100_1011001;
		logarithm_table[3323] = 14'b0000100_1011001;
		logarithm_table[3324] = 14'b0000100_1011001;
		logarithm_table[3325] = 14'b0000100_1011001;
		logarithm_table[3326] = 14'b0000100_1011010;
		logarithm_table[3327] = 14'b0000100_1011010;
		logarithm_table[3328] = 14'b0000100_1011010;
		logarithm_table[3329] = 14'b0000100_1011010;
		logarithm_table[3330] = 14'b0000100_1011010;
		logarithm_table[3331] = 14'b0000100_1011010;
		logarithm_table[3332] = 14'b0000100_1011010;
		logarithm_table[3333] = 14'b0000100_1011010;
		logarithm_table[3334] = 14'b0000100_1011010;
		logarithm_table[3335] = 14'b0000100_1011010;
		logarithm_table[3336] = 14'b0000100_1011010;
		logarithm_table[3337] = 14'b0000100_1011010;
		logarithm_table[3338] = 14'b0000100_1011010;
		logarithm_table[3339] = 14'b0000100_1011010;
		logarithm_table[3340] = 14'b0000100_1011010;
		logarithm_table[3341] = 14'b0000100_1011010;
		logarithm_table[3342] = 14'b0000100_1011010;
		logarithm_table[3343] = 14'b0000100_1011010;
		logarithm_table[3344] = 14'b0000100_1011011;
		logarithm_table[3345] = 14'b0000100_1011011;
		logarithm_table[3346] = 14'b0000100_1011011;
		logarithm_table[3347] = 14'b0000100_1011011;
		logarithm_table[3348] = 14'b0000100_1011011;
		logarithm_table[3349] = 14'b0000100_1011011;
		logarithm_table[3350] = 14'b0000100_1011011;
		logarithm_table[3351] = 14'b0000100_1011011;
		logarithm_table[3352] = 14'b0000100_1011011;
		logarithm_table[3353] = 14'b0000100_1011011;
		logarithm_table[3354] = 14'b0000100_1011011;
		logarithm_table[3355] = 14'b0000100_1011011;
		logarithm_table[3356] = 14'b0000100_1011011;
		logarithm_table[3357] = 14'b0000100_1011011;
		logarithm_table[3358] = 14'b0000100_1011011;
		logarithm_table[3359] = 14'b0000100_1011011;
		logarithm_table[3360] = 14'b0000100_1011011;
		logarithm_table[3361] = 14'b0000100_1011011;
		logarithm_table[3362] = 14'b0000100_1011100;
		logarithm_table[3363] = 14'b0000100_1011100;
		logarithm_table[3364] = 14'b0000100_1011100;
		logarithm_table[3365] = 14'b0000100_1011100;
		logarithm_table[3366] = 14'b0000100_1011100;
		logarithm_table[3367] = 14'b0000100_1011100;
		logarithm_table[3368] = 14'b0000100_1011100;
		logarithm_table[3369] = 14'b0000100_1011100;
		logarithm_table[3370] = 14'b0000100_1011100;
		logarithm_table[3371] = 14'b0000100_1011100;
		logarithm_table[3372] = 14'b0000100_1011100;
		logarithm_table[3373] = 14'b0000100_1011100;
		logarithm_table[3374] = 14'b0000100_1011100;
		logarithm_table[3375] = 14'b0000100_1011100;
		logarithm_table[3376] = 14'b0000100_1011100;
		logarithm_table[3377] = 14'b0000100_1011100;
		logarithm_table[3378] = 14'b0000100_1011100;
		logarithm_table[3379] = 14'b0000100_1011100;
		logarithm_table[3380] = 14'b0000100_1011101;
		logarithm_table[3381] = 14'b0000100_1011101;
		logarithm_table[3382] = 14'b0000100_1011101;
		logarithm_table[3383] = 14'b0000100_1011101;
		logarithm_table[3384] = 14'b0000100_1011101;
		logarithm_table[3385] = 14'b0000100_1011101;
		logarithm_table[3386] = 14'b0000100_1011101;
		logarithm_table[3387] = 14'b0000100_1011101;
		logarithm_table[3388] = 14'b0000100_1011101;
		logarithm_table[3389] = 14'b0000100_1011101;
		logarithm_table[3390] = 14'b0000100_1011101;
		logarithm_table[3391] = 14'b0000100_1011101;
		logarithm_table[3392] = 14'b0000100_1011101;
		logarithm_table[3393] = 14'b0000100_1011101;
		logarithm_table[3394] = 14'b0000100_1011101;
		logarithm_table[3395] = 14'b0000100_1011101;
		logarithm_table[3396] = 14'b0000100_1011101;
		logarithm_table[3397] = 14'b0000100_1011101;
		logarithm_table[3398] = 14'b0000100_1011110;
		logarithm_table[3399] = 14'b0000100_1011110;
		logarithm_table[3400] = 14'b0000100_1011110;
		logarithm_table[3401] = 14'b0000100_1011110;
		logarithm_table[3402] = 14'b0000100_1011110;
		logarithm_table[3403] = 14'b0000100_1011110;
		logarithm_table[3404] = 14'b0000100_1011110;
		logarithm_table[3405] = 14'b0000100_1011110;
		logarithm_table[3406] = 14'b0000100_1011110;
		logarithm_table[3407] = 14'b0000100_1011110;
		logarithm_table[3408] = 14'b0000100_1011110;
		logarithm_table[3409] = 14'b0000100_1011110;
		logarithm_table[3410] = 14'b0000100_1011110;
		logarithm_table[3411] = 14'b0000100_1011110;
		logarithm_table[3412] = 14'b0000100_1011110;
		logarithm_table[3413] = 14'b0000100_1011110;
		logarithm_table[3414] = 14'b0000100_1011110;
		logarithm_table[3415] = 14'b0000100_1011110;
		logarithm_table[3416] = 14'b0000100_1011110;
		logarithm_table[3417] = 14'b0000100_1011111;
		logarithm_table[3418] = 14'b0000100_1011111;
		logarithm_table[3419] = 14'b0000100_1011111;
		logarithm_table[3420] = 14'b0000100_1011111;
		logarithm_table[3421] = 14'b0000100_1011111;
		logarithm_table[3422] = 14'b0000100_1011111;
		logarithm_table[3423] = 14'b0000100_1011111;
		logarithm_table[3424] = 14'b0000100_1011111;
		logarithm_table[3425] = 14'b0000100_1011111;
		logarithm_table[3426] = 14'b0000100_1011111;
		logarithm_table[3427] = 14'b0000100_1011111;
		logarithm_table[3428] = 14'b0000100_1011111;
		logarithm_table[3429] = 14'b0000100_1011111;
		logarithm_table[3430] = 14'b0000100_1011111;
		logarithm_table[3431] = 14'b0000100_1011111;
		logarithm_table[3432] = 14'b0000100_1011111;
		logarithm_table[3433] = 14'b0000100_1011111;
		logarithm_table[3434] = 14'b0000100_1011111;
		logarithm_table[3435] = 14'b0000100_1100000;
		logarithm_table[3436] = 14'b0000100_1100000;
		logarithm_table[3437] = 14'b0000100_1100000;
		logarithm_table[3438] = 14'b0000100_1100000;
		logarithm_table[3439] = 14'b0000100_1100000;
		logarithm_table[3440] = 14'b0000100_1100000;
		logarithm_table[3441] = 14'b0000100_1100000;
		logarithm_table[3442] = 14'b0000100_1100000;
		logarithm_table[3443] = 14'b0000100_1100000;
		logarithm_table[3444] = 14'b0000100_1100000;
		logarithm_table[3445] = 14'b0000100_1100000;
		logarithm_table[3446] = 14'b0000100_1100000;
		logarithm_table[3447] = 14'b0000100_1100000;
		logarithm_table[3448] = 14'b0000100_1100000;
		logarithm_table[3449] = 14'b0000100_1100000;
		logarithm_table[3450] = 14'b0000100_1100000;
		logarithm_table[3451] = 14'b0000100_1100000;
		logarithm_table[3452] = 14'b0000100_1100000;
		logarithm_table[3453] = 14'b0000100_1100000;
		logarithm_table[3454] = 14'b0000100_1100001;
		logarithm_table[3455] = 14'b0000100_1100001;
		logarithm_table[3456] = 14'b0000100_1100001;
		logarithm_table[3457] = 14'b0000100_1100001;
		logarithm_table[3458] = 14'b0000100_1100001;
		logarithm_table[3459] = 14'b0000100_1100001;
		logarithm_table[3460] = 14'b0000100_1100001;
		logarithm_table[3461] = 14'b0000100_1100001;
		logarithm_table[3462] = 14'b0000100_1100001;
		logarithm_table[3463] = 14'b0000100_1100001;
		logarithm_table[3464] = 14'b0000100_1100001;
		logarithm_table[3465] = 14'b0000100_1100001;
		logarithm_table[3466] = 14'b0000100_1100001;
		logarithm_table[3467] = 14'b0000100_1100001;
		logarithm_table[3468] = 14'b0000100_1100001;
		logarithm_table[3469] = 14'b0000100_1100001;
		logarithm_table[3470] = 14'b0000100_1100001;
		logarithm_table[3471] = 14'b0000100_1100001;
		logarithm_table[3472] = 14'b0000100_1100001;
		logarithm_table[3473] = 14'b0000100_1100010;
		logarithm_table[3474] = 14'b0000100_1100010;
		logarithm_table[3475] = 14'b0000100_1100010;
		logarithm_table[3476] = 14'b0000100_1100010;
		logarithm_table[3477] = 14'b0000100_1100010;
		logarithm_table[3478] = 14'b0000100_1100010;
		logarithm_table[3479] = 14'b0000100_1100010;
		logarithm_table[3480] = 14'b0000100_1100010;
		logarithm_table[3481] = 14'b0000100_1100010;
		logarithm_table[3482] = 14'b0000100_1100010;
		logarithm_table[3483] = 14'b0000100_1100010;
		logarithm_table[3484] = 14'b0000100_1100010;
		logarithm_table[3485] = 14'b0000100_1100010;
		logarithm_table[3486] = 14'b0000100_1100010;
		logarithm_table[3487] = 14'b0000100_1100010;
		logarithm_table[3488] = 14'b0000100_1100010;
		logarithm_table[3489] = 14'b0000100_1100010;
		logarithm_table[3490] = 14'b0000100_1100010;
		logarithm_table[3491] = 14'b0000100_1100010;
		logarithm_table[3492] = 14'b0000100_1100011;
		logarithm_table[3493] = 14'b0000100_1100011;
		logarithm_table[3494] = 14'b0000100_1100011;
		logarithm_table[3495] = 14'b0000100_1100011;
		logarithm_table[3496] = 14'b0000100_1100011;
		logarithm_table[3497] = 14'b0000100_1100011;
		logarithm_table[3498] = 14'b0000100_1100011;
		logarithm_table[3499] = 14'b0000100_1100011;
		logarithm_table[3500] = 14'b0000100_1100011;
		logarithm_table[3501] = 14'b0000100_1100011;
		logarithm_table[3502] = 14'b0000100_1100011;
		logarithm_table[3503] = 14'b0000100_1100011;
		logarithm_table[3504] = 14'b0000100_1100011;
		logarithm_table[3505] = 14'b0000100_1100011;
		logarithm_table[3506] = 14'b0000100_1100011;
		logarithm_table[3507] = 14'b0000100_1100011;
		logarithm_table[3508] = 14'b0000100_1100011;
		logarithm_table[3509] = 14'b0000100_1100011;
		logarithm_table[3510] = 14'b0000100_1100011;
		logarithm_table[3511] = 14'b0000100_1100100;
		logarithm_table[3512] = 14'b0000100_1100100;
		logarithm_table[3513] = 14'b0000100_1100100;
		logarithm_table[3514] = 14'b0000100_1100100;
		logarithm_table[3515] = 14'b0000100_1100100;
		logarithm_table[3516] = 14'b0000100_1100100;
		logarithm_table[3517] = 14'b0000100_1100100;
		logarithm_table[3518] = 14'b0000100_1100100;
		logarithm_table[3519] = 14'b0000100_1100100;
		logarithm_table[3520] = 14'b0000100_1100100;
		logarithm_table[3521] = 14'b0000100_1100100;
		logarithm_table[3522] = 14'b0000100_1100100;
		logarithm_table[3523] = 14'b0000100_1100100;
		logarithm_table[3524] = 14'b0000100_1100100;
		logarithm_table[3525] = 14'b0000100_1100100;
		logarithm_table[3526] = 14'b0000100_1100100;
		logarithm_table[3527] = 14'b0000100_1100100;
		logarithm_table[3528] = 14'b0000100_1100100;
		logarithm_table[3529] = 14'b0000100_1100100;
		logarithm_table[3530] = 14'b0000100_1100101;
		logarithm_table[3531] = 14'b0000100_1100101;
		logarithm_table[3532] = 14'b0000100_1100101;
		logarithm_table[3533] = 14'b0000100_1100101;
		logarithm_table[3534] = 14'b0000100_1100101;
		logarithm_table[3535] = 14'b0000100_1100101;
		logarithm_table[3536] = 14'b0000100_1100101;
		logarithm_table[3537] = 14'b0000100_1100101;
		logarithm_table[3538] = 14'b0000100_1100101;
		logarithm_table[3539] = 14'b0000100_1100101;
		logarithm_table[3540] = 14'b0000100_1100101;
		logarithm_table[3541] = 14'b0000100_1100101;
		logarithm_table[3542] = 14'b0000100_1100101;
		logarithm_table[3543] = 14'b0000100_1100101;
		logarithm_table[3544] = 14'b0000100_1100101;
		logarithm_table[3545] = 14'b0000100_1100101;
		logarithm_table[3546] = 14'b0000100_1100101;
		logarithm_table[3547] = 14'b0000100_1100101;
		logarithm_table[3548] = 14'b0000100_1100101;
		logarithm_table[3549] = 14'b0000100_1100110;
		logarithm_table[3550] = 14'b0000100_1100110;
		logarithm_table[3551] = 14'b0000100_1100110;
		logarithm_table[3552] = 14'b0000100_1100110;
		logarithm_table[3553] = 14'b0000100_1100110;
		logarithm_table[3554] = 14'b0000100_1100110;
		logarithm_table[3555] = 14'b0000100_1100110;
		logarithm_table[3556] = 14'b0000100_1100110;
		logarithm_table[3557] = 14'b0000100_1100110;
		logarithm_table[3558] = 14'b0000100_1100110;
		logarithm_table[3559] = 14'b0000100_1100110;
		logarithm_table[3560] = 14'b0000100_1100110;
		logarithm_table[3561] = 14'b0000100_1100110;
		logarithm_table[3562] = 14'b0000100_1100110;
		logarithm_table[3563] = 14'b0000100_1100110;
		logarithm_table[3564] = 14'b0000100_1100110;
		logarithm_table[3565] = 14'b0000100_1100110;
		logarithm_table[3566] = 14'b0000100_1100110;
		logarithm_table[3567] = 14'b0000100_1100110;
		logarithm_table[3568] = 14'b0000100_1100111;
		logarithm_table[3569] = 14'b0000100_1100111;
		logarithm_table[3570] = 14'b0000100_1100111;
		logarithm_table[3571] = 14'b0000100_1100111;
		logarithm_table[3572] = 14'b0000100_1100111;
		logarithm_table[3573] = 14'b0000100_1100111;
		logarithm_table[3574] = 14'b0000100_1100111;
		logarithm_table[3575] = 14'b0000100_1100111;
		logarithm_table[3576] = 14'b0000100_1100111;
		logarithm_table[3577] = 14'b0000100_1100111;
		logarithm_table[3578] = 14'b0000100_1100111;
		logarithm_table[3579] = 14'b0000100_1100111;
		logarithm_table[3580] = 14'b0000100_1100111;
		logarithm_table[3581] = 14'b0000100_1100111;
		logarithm_table[3582] = 14'b0000100_1100111;
		logarithm_table[3583] = 14'b0000100_1100111;
		logarithm_table[3584] = 14'b0000100_1100111;
		logarithm_table[3585] = 14'b0000100_1100111;
		logarithm_table[3586] = 14'b0000100_1100111;
		logarithm_table[3587] = 14'b0000100_1100111;
		logarithm_table[3588] = 14'b0000100_1101000;
		logarithm_table[3589] = 14'b0000100_1101000;
		logarithm_table[3590] = 14'b0000100_1101000;
		logarithm_table[3591] = 14'b0000100_1101000;
		logarithm_table[3592] = 14'b0000100_1101000;
		logarithm_table[3593] = 14'b0000100_1101000;
		logarithm_table[3594] = 14'b0000100_1101000;
		logarithm_table[3595] = 14'b0000100_1101000;
		logarithm_table[3596] = 14'b0000100_1101000;
		logarithm_table[3597] = 14'b0000100_1101000;
		logarithm_table[3598] = 14'b0000100_1101000;
		logarithm_table[3599] = 14'b0000100_1101000;
		logarithm_table[3600] = 14'b0000100_1101000;
		logarithm_table[3601] = 14'b0000100_1101000;
		logarithm_table[3602] = 14'b0000100_1101000;
		logarithm_table[3603] = 14'b0000100_1101000;
		logarithm_table[3604] = 14'b0000100_1101000;
		logarithm_table[3605] = 14'b0000100_1101000;
		logarithm_table[3606] = 14'b0000100_1101000;
		logarithm_table[3607] = 14'b0000100_1101001;
		logarithm_table[3608] = 14'b0000100_1101001;
		logarithm_table[3609] = 14'b0000100_1101001;
		logarithm_table[3610] = 14'b0000100_1101001;
		logarithm_table[3611] = 14'b0000100_1101001;
		logarithm_table[3612] = 14'b0000100_1101001;
		logarithm_table[3613] = 14'b0000100_1101001;
		logarithm_table[3614] = 14'b0000100_1101001;
		logarithm_table[3615] = 14'b0000100_1101001;
		logarithm_table[3616] = 14'b0000100_1101001;
		logarithm_table[3617] = 14'b0000100_1101001;
		logarithm_table[3618] = 14'b0000100_1101001;
		logarithm_table[3619] = 14'b0000100_1101001;
		logarithm_table[3620] = 14'b0000100_1101001;
		logarithm_table[3621] = 14'b0000100_1101001;
		logarithm_table[3622] = 14'b0000100_1101001;
		logarithm_table[3623] = 14'b0000100_1101001;
		logarithm_table[3624] = 14'b0000100_1101001;
		logarithm_table[3625] = 14'b0000100_1101001;
		logarithm_table[3626] = 14'b0000100_1101001;
		logarithm_table[3627] = 14'b0000100_1101010;
		logarithm_table[3628] = 14'b0000100_1101010;
		logarithm_table[3629] = 14'b0000100_1101010;
		logarithm_table[3630] = 14'b0000100_1101010;
		logarithm_table[3631] = 14'b0000100_1101010;
		logarithm_table[3632] = 14'b0000100_1101010;
		logarithm_table[3633] = 14'b0000100_1101010;
		logarithm_table[3634] = 14'b0000100_1101010;
		logarithm_table[3635] = 14'b0000100_1101010;
		logarithm_table[3636] = 14'b0000100_1101010;
		logarithm_table[3637] = 14'b0000100_1101010;
		logarithm_table[3638] = 14'b0000100_1101010;
		logarithm_table[3639] = 14'b0000100_1101010;
		logarithm_table[3640] = 14'b0000100_1101010;
		logarithm_table[3641] = 14'b0000100_1101010;
		logarithm_table[3642] = 14'b0000100_1101010;
		logarithm_table[3643] = 14'b0000100_1101010;
		logarithm_table[3644] = 14'b0000100_1101010;
		logarithm_table[3645] = 14'b0000100_1101010;
		logarithm_table[3646] = 14'b0000100_1101011;
		logarithm_table[3647] = 14'b0000100_1101011;
		logarithm_table[3648] = 14'b0000100_1101011;
		logarithm_table[3649] = 14'b0000100_1101011;
		logarithm_table[3650] = 14'b0000100_1101011;
		logarithm_table[3651] = 14'b0000100_1101011;
		logarithm_table[3652] = 14'b0000100_1101011;
		logarithm_table[3653] = 14'b0000100_1101011;
		logarithm_table[3654] = 14'b0000100_1101011;
		logarithm_table[3655] = 14'b0000100_1101011;
		logarithm_table[3656] = 14'b0000100_1101011;
		logarithm_table[3657] = 14'b0000100_1101011;
		logarithm_table[3658] = 14'b0000100_1101011;
		logarithm_table[3659] = 14'b0000100_1101011;
		logarithm_table[3660] = 14'b0000100_1101011;
		logarithm_table[3661] = 14'b0000100_1101011;
		logarithm_table[3662] = 14'b0000100_1101011;
		logarithm_table[3663] = 14'b0000100_1101011;
		logarithm_table[3664] = 14'b0000100_1101011;
		logarithm_table[3665] = 14'b0000100_1101011;
		logarithm_table[3666] = 14'b0000100_1101100;
		logarithm_table[3667] = 14'b0000100_1101100;
		logarithm_table[3668] = 14'b0000100_1101100;
		logarithm_table[3669] = 14'b0000100_1101100;
		logarithm_table[3670] = 14'b0000100_1101100;
		logarithm_table[3671] = 14'b0000100_1101100;
		logarithm_table[3672] = 14'b0000100_1101100;
		logarithm_table[3673] = 14'b0000100_1101100;
		logarithm_table[3674] = 14'b0000100_1101100;
		logarithm_table[3675] = 14'b0000100_1101100;
		logarithm_table[3676] = 14'b0000100_1101100;
		logarithm_table[3677] = 14'b0000100_1101100;
		logarithm_table[3678] = 14'b0000100_1101100;
		logarithm_table[3679] = 14'b0000100_1101100;
		logarithm_table[3680] = 14'b0000100_1101100;
		logarithm_table[3681] = 14'b0000100_1101100;
		logarithm_table[3682] = 14'b0000100_1101100;
		logarithm_table[3683] = 14'b0000100_1101100;
		logarithm_table[3684] = 14'b0000100_1101100;
		logarithm_table[3685] = 14'b0000100_1101100;
		logarithm_table[3686] = 14'b0000100_1101101;
		logarithm_table[3687] = 14'b0000100_1101101;
		logarithm_table[3688] = 14'b0000100_1101101;
		logarithm_table[3689] = 14'b0000100_1101101;
		logarithm_table[3690] = 14'b0000100_1101101;
		logarithm_table[3691] = 14'b0000100_1101101;
		logarithm_table[3692] = 14'b0000100_1101101;
		logarithm_table[3693] = 14'b0000100_1101101;
		logarithm_table[3694] = 14'b0000100_1101101;
		logarithm_table[3695] = 14'b0000100_1101101;
		logarithm_table[3696] = 14'b0000100_1101101;
		logarithm_table[3697] = 14'b0000100_1101101;
		logarithm_table[3698] = 14'b0000100_1101101;
		logarithm_table[3699] = 14'b0000100_1101101;
		logarithm_table[3700] = 14'b0000100_1101101;
		logarithm_table[3701] = 14'b0000100_1101101;
		logarithm_table[3702] = 14'b0000100_1101101;
		logarithm_table[3703] = 14'b0000100_1101101;
		logarithm_table[3704] = 14'b0000100_1101101;
		logarithm_table[3705] = 14'b0000100_1101101;
		logarithm_table[3706] = 14'b0000100_1101110;
		logarithm_table[3707] = 14'b0000100_1101110;
		logarithm_table[3708] = 14'b0000100_1101110;
		logarithm_table[3709] = 14'b0000100_1101110;
		logarithm_table[3710] = 14'b0000100_1101110;
		logarithm_table[3711] = 14'b0000100_1101110;
		logarithm_table[3712] = 14'b0000100_1101110;
		logarithm_table[3713] = 14'b0000100_1101110;
		logarithm_table[3714] = 14'b0000100_1101110;
		logarithm_table[3715] = 14'b0000100_1101110;
		logarithm_table[3716] = 14'b0000100_1101110;
		logarithm_table[3717] = 14'b0000100_1101110;
		logarithm_table[3718] = 14'b0000100_1101110;
		logarithm_table[3719] = 14'b0000100_1101110;
		logarithm_table[3720] = 14'b0000100_1101110;
		logarithm_table[3721] = 14'b0000100_1101110;
		logarithm_table[3722] = 14'b0000100_1101110;
		logarithm_table[3723] = 14'b0000100_1101110;
		logarithm_table[3724] = 14'b0000100_1101110;
		logarithm_table[3725] = 14'b0000100_1101110;
		logarithm_table[3726] = 14'b0000100_1101111;
		logarithm_table[3727] = 14'b0000100_1101111;
		logarithm_table[3728] = 14'b0000100_1101111;
		logarithm_table[3729] = 14'b0000100_1101111;
		logarithm_table[3730] = 14'b0000100_1101111;
		logarithm_table[3731] = 14'b0000100_1101111;
		logarithm_table[3732] = 14'b0000100_1101111;
		logarithm_table[3733] = 14'b0000100_1101111;
		logarithm_table[3734] = 14'b0000100_1101111;
		logarithm_table[3735] = 14'b0000100_1101111;
		logarithm_table[3736] = 14'b0000100_1101111;
		logarithm_table[3737] = 14'b0000100_1101111;
		logarithm_table[3738] = 14'b0000100_1101111;
		logarithm_table[3739] = 14'b0000100_1101111;
		logarithm_table[3740] = 14'b0000100_1101111;
		logarithm_table[3741] = 14'b0000100_1101111;
		logarithm_table[3742] = 14'b0000100_1101111;
		logarithm_table[3743] = 14'b0000100_1101111;
		logarithm_table[3744] = 14'b0000100_1101111;
		logarithm_table[3745] = 14'b0000100_1101111;
		logarithm_table[3746] = 14'b0000100_1110000;
		logarithm_table[3747] = 14'b0000100_1110000;
		logarithm_table[3748] = 14'b0000100_1110000;
		logarithm_table[3749] = 14'b0000100_1110000;
		logarithm_table[3750] = 14'b0000100_1110000;
		logarithm_table[3751] = 14'b0000100_1110000;
		logarithm_table[3752] = 14'b0000100_1110000;
		logarithm_table[3753] = 14'b0000100_1110000;
		logarithm_table[3754] = 14'b0000100_1110000;
		logarithm_table[3755] = 14'b0000100_1110000;
		logarithm_table[3756] = 14'b0000100_1110000;
		logarithm_table[3757] = 14'b0000100_1110000;
		logarithm_table[3758] = 14'b0000100_1110000;
		logarithm_table[3759] = 14'b0000100_1110000;
		logarithm_table[3760] = 14'b0000100_1110000;
		logarithm_table[3761] = 14'b0000100_1110000;
		logarithm_table[3762] = 14'b0000100_1110000;
		logarithm_table[3763] = 14'b0000100_1110000;
		logarithm_table[3764] = 14'b0000100_1110000;
		logarithm_table[3765] = 14'b0000100_1110000;
		logarithm_table[3766] = 14'b0000100_1110000;
		logarithm_table[3767] = 14'b0000100_1110001;
		logarithm_table[3768] = 14'b0000100_1110001;
		logarithm_table[3769] = 14'b0000100_1110001;
		logarithm_table[3770] = 14'b0000100_1110001;
		logarithm_table[3771] = 14'b0000100_1110001;
		logarithm_table[3772] = 14'b0000100_1110001;
		logarithm_table[3773] = 14'b0000100_1110001;
		logarithm_table[3774] = 14'b0000100_1110001;
		logarithm_table[3775] = 14'b0000100_1110001;
		logarithm_table[3776] = 14'b0000100_1110001;
		logarithm_table[3777] = 14'b0000100_1110001;
		logarithm_table[3778] = 14'b0000100_1110001;
		logarithm_table[3779] = 14'b0000100_1110001;
		logarithm_table[3780] = 14'b0000100_1110001;
		logarithm_table[3781] = 14'b0000100_1110001;
		logarithm_table[3782] = 14'b0000100_1110001;
		logarithm_table[3783] = 14'b0000100_1110001;
		logarithm_table[3784] = 14'b0000100_1110001;
		logarithm_table[3785] = 14'b0000100_1110001;
		logarithm_table[3786] = 14'b0000100_1110001;
		logarithm_table[3787] = 14'b0000100_1110010;
		logarithm_table[3788] = 14'b0000100_1110010;
		logarithm_table[3789] = 14'b0000100_1110010;
		logarithm_table[3790] = 14'b0000100_1110010;
		logarithm_table[3791] = 14'b0000100_1110010;
		logarithm_table[3792] = 14'b0000100_1110010;
		logarithm_table[3793] = 14'b0000100_1110010;
		logarithm_table[3794] = 14'b0000100_1110010;
		logarithm_table[3795] = 14'b0000100_1110010;
		logarithm_table[3796] = 14'b0000100_1110010;
		logarithm_table[3797] = 14'b0000100_1110010;
		logarithm_table[3798] = 14'b0000100_1110010;
		logarithm_table[3799] = 14'b0000100_1110010;
		logarithm_table[3800] = 14'b0000100_1110010;
		logarithm_table[3801] = 14'b0000100_1110010;
		logarithm_table[3802] = 14'b0000100_1110010;
		logarithm_table[3803] = 14'b0000100_1110010;
		logarithm_table[3804] = 14'b0000100_1110010;
		logarithm_table[3805] = 14'b0000100_1110010;
		logarithm_table[3806] = 14'b0000100_1110010;
		logarithm_table[3807] = 14'b0000100_1110010;
		logarithm_table[3808] = 14'b0000100_1110011;
		logarithm_table[3809] = 14'b0000100_1110011;
		logarithm_table[3810] = 14'b0000100_1110011;
		logarithm_table[3811] = 14'b0000100_1110011;
		logarithm_table[3812] = 14'b0000100_1110011;
		logarithm_table[3813] = 14'b0000100_1110011;
		logarithm_table[3814] = 14'b0000100_1110011;
		logarithm_table[3815] = 14'b0000100_1110011;
		logarithm_table[3816] = 14'b0000100_1110011;
		logarithm_table[3817] = 14'b0000100_1110011;
		logarithm_table[3818] = 14'b0000100_1110011;
		logarithm_table[3819] = 14'b0000100_1110011;
		logarithm_table[3820] = 14'b0000100_1110011;
		logarithm_table[3821] = 14'b0000100_1110011;
		logarithm_table[3822] = 14'b0000100_1110011;
		logarithm_table[3823] = 14'b0000100_1110011;
		logarithm_table[3824] = 14'b0000100_1110011;
		logarithm_table[3825] = 14'b0000100_1110011;
		logarithm_table[3826] = 14'b0000100_1110011;
		logarithm_table[3827] = 14'b0000100_1110011;
		logarithm_table[3828] = 14'b0000100_1110100;
		logarithm_table[3829] = 14'b0000100_1110100;
		logarithm_table[3830] = 14'b0000100_1110100;
		logarithm_table[3831] = 14'b0000100_1110100;
		logarithm_table[3832] = 14'b0000100_1110100;
		logarithm_table[3833] = 14'b0000100_1110100;
		logarithm_table[3834] = 14'b0000100_1110100;
		logarithm_table[3835] = 14'b0000100_1110100;
		logarithm_table[3836] = 14'b0000100_1110100;
		logarithm_table[3837] = 14'b0000100_1110100;
		logarithm_table[3838] = 14'b0000100_1110100;
		logarithm_table[3839] = 14'b0000100_1110100;
		logarithm_table[3840] = 14'b0000100_1110100;
		logarithm_table[3841] = 14'b0000100_1110100;
		logarithm_table[3842] = 14'b0000100_1110100;
		logarithm_table[3843] = 14'b0000100_1110100;
		logarithm_table[3844] = 14'b0000100_1110100;
		logarithm_table[3845] = 14'b0000100_1110100;
		logarithm_table[3846] = 14'b0000100_1110100;
		logarithm_table[3847] = 14'b0000100_1110100;
		logarithm_table[3848] = 14'b0000100_1110100;
		logarithm_table[3849] = 14'b0000100_1110101;
		logarithm_table[3850] = 14'b0000100_1110101;
		logarithm_table[3851] = 14'b0000100_1110101;
		logarithm_table[3852] = 14'b0000100_1110101;
		logarithm_table[3853] = 14'b0000100_1110101;
		logarithm_table[3854] = 14'b0000100_1110101;
		logarithm_table[3855] = 14'b0000100_1110101;
		logarithm_table[3856] = 14'b0000100_1110101;
		logarithm_table[3857] = 14'b0000100_1110101;
		logarithm_table[3858] = 14'b0000100_1110101;
		logarithm_table[3859] = 14'b0000100_1110101;
		logarithm_table[3860] = 14'b0000100_1110101;
		logarithm_table[3861] = 14'b0000100_1110101;
		logarithm_table[3862] = 14'b0000100_1110101;
		logarithm_table[3863] = 14'b0000100_1110101;
		logarithm_table[3864] = 14'b0000100_1110101;
		logarithm_table[3865] = 14'b0000100_1110101;
		logarithm_table[3866] = 14'b0000100_1110101;
		logarithm_table[3867] = 14'b0000100_1110101;
		logarithm_table[3868] = 14'b0000100_1110101;
		logarithm_table[3869] = 14'b0000100_1110101;
		logarithm_table[3870] = 14'b0000100_1110110;
		logarithm_table[3871] = 14'b0000100_1110110;
		logarithm_table[3872] = 14'b0000100_1110110;
		logarithm_table[3873] = 14'b0000100_1110110;
		logarithm_table[3874] = 14'b0000100_1110110;
		logarithm_table[3875] = 14'b0000100_1110110;
		logarithm_table[3876] = 14'b0000100_1110110;
		logarithm_table[3877] = 14'b0000100_1110110;
		logarithm_table[3878] = 14'b0000100_1110110;
		logarithm_table[3879] = 14'b0000100_1110110;
		logarithm_table[3880] = 14'b0000100_1110110;
		logarithm_table[3881] = 14'b0000100_1110110;
		logarithm_table[3882] = 14'b0000100_1110110;
		logarithm_table[3883] = 14'b0000100_1110110;
		logarithm_table[3884] = 14'b0000100_1110110;
		logarithm_table[3885] = 14'b0000100_1110110;
		logarithm_table[3886] = 14'b0000100_1110110;
		logarithm_table[3887] = 14'b0000100_1110110;
		logarithm_table[3888] = 14'b0000100_1110110;
		logarithm_table[3889] = 14'b0000100_1110110;
		logarithm_table[3890] = 14'b0000100_1110110;
		logarithm_table[3891] = 14'b0000100_1110111;
		logarithm_table[3892] = 14'b0000100_1110111;
		logarithm_table[3893] = 14'b0000100_1110111;
		logarithm_table[3894] = 14'b0000100_1110111;
		logarithm_table[3895] = 14'b0000100_1110111;
		logarithm_table[3896] = 14'b0000100_1110111;
		logarithm_table[3897] = 14'b0000100_1110111;
		logarithm_table[3898] = 14'b0000100_1110111;
		logarithm_table[3899] = 14'b0000100_1110111;
		logarithm_table[3900] = 14'b0000100_1110111;
		logarithm_table[3901] = 14'b0000100_1110111;
		logarithm_table[3902] = 14'b0000100_1110111;
		logarithm_table[3903] = 14'b0000100_1110111;
		logarithm_table[3904] = 14'b0000100_1110111;
		logarithm_table[3905] = 14'b0000100_1110111;
		logarithm_table[3906] = 14'b0000100_1110111;
		logarithm_table[3907] = 14'b0000100_1110111;
		logarithm_table[3908] = 14'b0000100_1110111;
		logarithm_table[3909] = 14'b0000100_1110111;
		logarithm_table[3910] = 14'b0000100_1110111;
		logarithm_table[3911] = 14'b0000100_1110111;
		logarithm_table[3912] = 14'b0000100_1111000;
		logarithm_table[3913] = 14'b0000100_1111000;
		logarithm_table[3914] = 14'b0000100_1111000;
		logarithm_table[3915] = 14'b0000100_1111000;
		logarithm_table[3916] = 14'b0000100_1111000;
		logarithm_table[3917] = 14'b0000100_1111000;
		logarithm_table[3918] = 14'b0000100_1111000;
		logarithm_table[3919] = 14'b0000100_1111000;
		logarithm_table[3920] = 14'b0000100_1111000;
		logarithm_table[3921] = 14'b0000100_1111000;
		logarithm_table[3922] = 14'b0000100_1111000;
		logarithm_table[3923] = 14'b0000100_1111000;
		logarithm_table[3924] = 14'b0000100_1111000;
		logarithm_table[3925] = 14'b0000100_1111000;
		logarithm_table[3926] = 14'b0000100_1111000;
		logarithm_table[3927] = 14'b0000100_1111000;
		logarithm_table[3928] = 14'b0000100_1111000;
		logarithm_table[3929] = 14'b0000100_1111000;
		logarithm_table[3930] = 14'b0000100_1111000;
		logarithm_table[3931] = 14'b0000100_1111000;
		logarithm_table[3932] = 14'b0000100_1111000;
		logarithm_table[3933] = 14'b0000100_1111001;
		logarithm_table[3934] = 14'b0000100_1111001;
		logarithm_table[3935] = 14'b0000100_1111001;
		logarithm_table[3936] = 14'b0000100_1111001;
		logarithm_table[3937] = 14'b0000100_1111001;
		logarithm_table[3938] = 14'b0000100_1111001;
		logarithm_table[3939] = 14'b0000100_1111001;
		logarithm_table[3940] = 14'b0000100_1111001;
		logarithm_table[3941] = 14'b0000100_1111001;
		logarithm_table[3942] = 14'b0000100_1111001;
		logarithm_table[3943] = 14'b0000100_1111001;
		logarithm_table[3944] = 14'b0000100_1111001;
		logarithm_table[3945] = 14'b0000100_1111001;
		logarithm_table[3946] = 14'b0000100_1111001;
		logarithm_table[3947] = 14'b0000100_1111001;
		logarithm_table[3948] = 14'b0000100_1111001;
		logarithm_table[3949] = 14'b0000100_1111001;
		logarithm_table[3950] = 14'b0000100_1111001;
		logarithm_table[3951] = 14'b0000100_1111001;
		logarithm_table[3952] = 14'b0000100_1111001;
		logarithm_table[3953] = 14'b0000100_1111001;
		logarithm_table[3954] = 14'b0000100_1111001;
		logarithm_table[3955] = 14'b0000100_1111010;
		logarithm_table[3956] = 14'b0000100_1111010;
		logarithm_table[3957] = 14'b0000100_1111010;
		logarithm_table[3958] = 14'b0000100_1111010;
		logarithm_table[3959] = 14'b0000100_1111010;
		logarithm_table[3960] = 14'b0000100_1111010;
		logarithm_table[3961] = 14'b0000100_1111010;
		logarithm_table[3962] = 14'b0000100_1111010;
		logarithm_table[3963] = 14'b0000100_1111010;
		logarithm_table[3964] = 14'b0000100_1111010;
		logarithm_table[3965] = 14'b0000100_1111010;
		logarithm_table[3966] = 14'b0000100_1111010;
		logarithm_table[3967] = 14'b0000100_1111010;
		logarithm_table[3968] = 14'b0000100_1111010;
		logarithm_table[3969] = 14'b0000100_1111010;
		logarithm_table[3970] = 14'b0000100_1111010;
		logarithm_table[3971] = 14'b0000100_1111010;
		logarithm_table[3972] = 14'b0000100_1111010;
		logarithm_table[3973] = 14'b0000100_1111010;
		logarithm_table[3974] = 14'b0000100_1111010;
		logarithm_table[3975] = 14'b0000100_1111010;
		logarithm_table[3976] = 14'b0000100_1111011;
		logarithm_table[3977] = 14'b0000100_1111011;
		logarithm_table[3978] = 14'b0000100_1111011;
		logarithm_table[3979] = 14'b0000100_1111011;
		logarithm_table[3980] = 14'b0000100_1111011;
		logarithm_table[3981] = 14'b0000100_1111011;
		logarithm_table[3982] = 14'b0000100_1111011;
		logarithm_table[3983] = 14'b0000100_1111011;
		logarithm_table[3984] = 14'b0000100_1111011;
		logarithm_table[3985] = 14'b0000100_1111011;
		logarithm_table[3986] = 14'b0000100_1111011;
		logarithm_table[3987] = 14'b0000100_1111011;
		logarithm_table[3988] = 14'b0000100_1111011;
		logarithm_table[3989] = 14'b0000100_1111011;
		logarithm_table[3990] = 14'b0000100_1111011;
		logarithm_table[3991] = 14'b0000100_1111011;
		logarithm_table[3992] = 14'b0000100_1111011;
		logarithm_table[3993] = 14'b0000100_1111011;
		logarithm_table[3994] = 14'b0000100_1111011;
		logarithm_table[3995] = 14'b0000100_1111011;
		logarithm_table[3996] = 14'b0000100_1111011;
		logarithm_table[3997] = 14'b0000100_1111011;
		logarithm_table[3998] = 14'b0000100_1111100;
		logarithm_table[3999] = 14'b0000100_1111100;
		logarithm_table[4000] = 14'b0000100_1111100;
		logarithm_table[4001] = 14'b0000100_1111100;
		logarithm_table[4002] = 14'b0000100_1111100;
		logarithm_table[4003] = 14'b0000100_1111100;
		logarithm_table[4004] = 14'b0000100_1111100;
		logarithm_table[4005] = 14'b0000100_1111100;
		logarithm_table[4006] = 14'b0000100_1111100;
		logarithm_table[4007] = 14'b0000100_1111100;
		logarithm_table[4008] = 14'b0000100_1111100;
		logarithm_table[4009] = 14'b0000100_1111100;
		logarithm_table[4010] = 14'b0000100_1111100;
		logarithm_table[4011] = 14'b0000100_1111100;
		logarithm_table[4012] = 14'b0000100_1111100;
		logarithm_table[4013] = 14'b0000100_1111100;
		logarithm_table[4014] = 14'b0000100_1111100;
		logarithm_table[4015] = 14'b0000100_1111100;
		logarithm_table[4016] = 14'b0000100_1111100;
		logarithm_table[4017] = 14'b0000100_1111100;
		logarithm_table[4018] = 14'b0000100_1111100;
		logarithm_table[4019] = 14'b0000100_1111100;
		logarithm_table[4020] = 14'b0000100_1111101;
		logarithm_table[4021] = 14'b0000100_1111101;
		logarithm_table[4022] = 14'b0000100_1111101;
		logarithm_table[4023] = 14'b0000100_1111101;
		logarithm_table[4024] = 14'b0000100_1111101;
		logarithm_table[4025] = 14'b0000100_1111101;
		logarithm_table[4026] = 14'b0000100_1111101;
		logarithm_table[4027] = 14'b0000100_1111101;
		logarithm_table[4028] = 14'b0000100_1111101;
		logarithm_table[4029] = 14'b0000100_1111101;
		logarithm_table[4030] = 14'b0000100_1111101;
		logarithm_table[4031] = 14'b0000100_1111101;
		logarithm_table[4032] = 14'b0000100_1111101;
		logarithm_table[4033] = 14'b0000100_1111101;
		logarithm_table[4034] = 14'b0000100_1111101;
		logarithm_table[4035] = 14'b0000100_1111101;
		logarithm_table[4036] = 14'b0000100_1111101;
		logarithm_table[4037] = 14'b0000100_1111101;
		logarithm_table[4038] = 14'b0000100_1111101;
		logarithm_table[4039] = 14'b0000100_1111101;
		logarithm_table[4040] = 14'b0000100_1111101;
		logarithm_table[4041] = 14'b0000100_1111110;
		logarithm_table[4042] = 14'b0000100_1111110;
		logarithm_table[4043] = 14'b0000100_1111110;
		logarithm_table[4044] = 14'b0000100_1111110;
		logarithm_table[4045] = 14'b0000100_1111110;
		logarithm_table[4046] = 14'b0000100_1111110;
		logarithm_table[4047] = 14'b0000100_1111110;
		logarithm_table[4048] = 14'b0000100_1111110;
		logarithm_table[4049] = 14'b0000100_1111110;
		logarithm_table[4050] = 14'b0000100_1111110;
		logarithm_table[4051] = 14'b0000100_1111110;
		logarithm_table[4052] = 14'b0000100_1111110;
		logarithm_table[4053] = 14'b0000100_1111110;
		logarithm_table[4054] = 14'b0000100_1111110;
		logarithm_table[4055] = 14'b0000100_1111110;
		logarithm_table[4056] = 14'b0000100_1111110;
		logarithm_table[4057] = 14'b0000100_1111110;
		logarithm_table[4058] = 14'b0000100_1111110;
		logarithm_table[4059] = 14'b0000100_1111110;
		logarithm_table[4060] = 14'b0000100_1111110;
		logarithm_table[4061] = 14'b0000100_1111110;
		logarithm_table[4062] = 14'b0000100_1111110;
		logarithm_table[4063] = 14'b0000100_1111111;
		logarithm_table[4064] = 14'b0000100_1111111;
		logarithm_table[4065] = 14'b0000100_1111111;
		logarithm_table[4066] = 14'b0000100_1111111;
		logarithm_table[4067] = 14'b0000100_1111111;
		logarithm_table[4068] = 14'b0000100_1111111;
		logarithm_table[4069] = 14'b0000100_1111111;
		logarithm_table[4070] = 14'b0000100_1111111;
		logarithm_table[4071] = 14'b0000100_1111111;
		logarithm_table[4072] = 14'b0000100_1111111;
		logarithm_table[4073] = 14'b0000100_1111111;
		logarithm_table[4074] = 14'b0000100_1111111;
		logarithm_table[4075] = 14'b0000100_1111111;
		logarithm_table[4076] = 14'b0000100_1111111;
		logarithm_table[4077] = 14'b0000100_1111111;
		logarithm_table[4078] = 14'b0000100_1111111;
		logarithm_table[4079] = 14'b0000100_1111111;
		logarithm_table[4080] = 14'b0000100_1111111;
		logarithm_table[4081] = 14'b0000100_1111111;
		logarithm_table[4082] = 14'b0000100_1111111;
		logarithm_table[4083] = 14'b0000100_1111111;
		logarithm_table[4084] = 14'b0000100_1111111;
		logarithm_table[4085] = 14'b0000101_0000000;
		logarithm_table[4086] = 14'b0000101_0000000;
		logarithm_table[4087] = 14'b0000101_0000000;
		logarithm_table[4088] = 14'b0000101_0000000;
		logarithm_table[4089] = 14'b0000101_0000000;
		logarithm_table[4090] = 14'b0000101_0000000;
		logarithm_table[4091] = 14'b0000101_0000000;
		logarithm_table[4092] = 14'b0000101_0000000;
		logarithm_table[4093] = 14'b0000101_0000000;
		logarithm_table[4094] = 14'b0000101_0000000;
		logarithm_table[4095] = 14'b0000101_0000000;
		logarithm_table[4096] = 14'b0000101_0000000;
		logarithm_table[4097] = 14'b0000101_0000000;
		logarithm_table[4098] = 14'b0000101_0000000;
		logarithm_table[4099] = 14'b0000101_0000000;
		logarithm_table[4100] = 14'b0000101_0000000;
		logarithm_table[4101] = 14'b0000101_0000000;
		logarithm_table[4102] = 14'b0000101_0000000;
		logarithm_table[4103] = 14'b0000101_0000000;
		logarithm_table[4104] = 14'b0000101_0000000;
		logarithm_table[4105] = 14'b0000101_0000000;
		logarithm_table[4106] = 14'b0000101_0000000;
		logarithm_table[4107] = 14'b0000101_0000000;
		logarithm_table[4108] = 14'b0000101_0000001;
		logarithm_table[4109] = 14'b0000101_0000001;
		logarithm_table[4110] = 14'b0000101_0000001;
		logarithm_table[4111] = 14'b0000101_0000001;
		logarithm_table[4112] = 14'b0000101_0000001;
		logarithm_table[4113] = 14'b0000101_0000001;
		logarithm_table[4114] = 14'b0000101_0000001;
		logarithm_table[4115] = 14'b0000101_0000001;
		logarithm_table[4116] = 14'b0000101_0000001;
		logarithm_table[4117] = 14'b0000101_0000001;
		logarithm_table[4118] = 14'b0000101_0000001;
		logarithm_table[4119] = 14'b0000101_0000001;
		logarithm_table[4120] = 14'b0000101_0000001;
		logarithm_table[4121] = 14'b0000101_0000001;
		logarithm_table[4122] = 14'b0000101_0000001;
		logarithm_table[4123] = 14'b0000101_0000001;
		logarithm_table[4124] = 14'b0000101_0000001;
		logarithm_table[4125] = 14'b0000101_0000001;
		logarithm_table[4126] = 14'b0000101_0000001;
		logarithm_table[4127] = 14'b0000101_0000001;
		logarithm_table[4128] = 14'b0000101_0000001;
		logarithm_table[4129] = 14'b0000101_0000001;
		logarithm_table[4130] = 14'b0000101_0000010;
		logarithm_table[4131] = 14'b0000101_0000010;
		logarithm_table[4132] = 14'b0000101_0000010;
		logarithm_table[4133] = 14'b0000101_0000010;
		logarithm_table[4134] = 14'b0000101_0000010;
		logarithm_table[4135] = 14'b0000101_0000010;
		logarithm_table[4136] = 14'b0000101_0000010;
		logarithm_table[4137] = 14'b0000101_0000010;
		logarithm_table[4138] = 14'b0000101_0000010;
		logarithm_table[4139] = 14'b0000101_0000010;
		logarithm_table[4140] = 14'b0000101_0000010;
		logarithm_table[4141] = 14'b0000101_0000010;
		logarithm_table[4142] = 14'b0000101_0000010;
		logarithm_table[4143] = 14'b0000101_0000010;
		logarithm_table[4144] = 14'b0000101_0000010;
		logarithm_table[4145] = 14'b0000101_0000010;
		logarithm_table[4146] = 14'b0000101_0000010;
		logarithm_table[4147] = 14'b0000101_0000010;
		logarithm_table[4148] = 14'b0000101_0000010;
		logarithm_table[4149] = 14'b0000101_0000010;
		logarithm_table[4150] = 14'b0000101_0000010;
		logarithm_table[4151] = 14'b0000101_0000010;
		logarithm_table[4152] = 14'b0000101_0000011;
		logarithm_table[4153] = 14'b0000101_0000011;
		logarithm_table[4154] = 14'b0000101_0000011;
		logarithm_table[4155] = 14'b0000101_0000011;
		logarithm_table[4156] = 14'b0000101_0000011;
		logarithm_table[4157] = 14'b0000101_0000011;
		logarithm_table[4158] = 14'b0000101_0000011;
		logarithm_table[4159] = 14'b0000101_0000011;
		logarithm_table[4160] = 14'b0000101_0000011;
		logarithm_table[4161] = 14'b0000101_0000011;
		logarithm_table[4162] = 14'b0000101_0000011;
		logarithm_table[4163] = 14'b0000101_0000011;
		logarithm_table[4164] = 14'b0000101_0000011;
		logarithm_table[4165] = 14'b0000101_0000011;
		logarithm_table[4166] = 14'b0000101_0000011;
		logarithm_table[4167] = 14'b0000101_0000011;
		logarithm_table[4168] = 14'b0000101_0000011;
		logarithm_table[4169] = 14'b0000101_0000011;
		logarithm_table[4170] = 14'b0000101_0000011;
		logarithm_table[4171] = 14'b0000101_0000011;
		logarithm_table[4172] = 14'b0000101_0000011;
		logarithm_table[4173] = 14'b0000101_0000011;
		logarithm_table[4174] = 14'b0000101_0000011;
		logarithm_table[4175] = 14'b0000101_0000100;
		logarithm_table[4176] = 14'b0000101_0000100;
		logarithm_table[4177] = 14'b0000101_0000100;
		logarithm_table[4178] = 14'b0000101_0000100;
		logarithm_table[4179] = 14'b0000101_0000100;
		logarithm_table[4180] = 14'b0000101_0000100;
		logarithm_table[4181] = 14'b0000101_0000100;
		logarithm_table[4182] = 14'b0000101_0000100;
		logarithm_table[4183] = 14'b0000101_0000100;
		logarithm_table[4184] = 14'b0000101_0000100;
		logarithm_table[4185] = 14'b0000101_0000100;
		logarithm_table[4186] = 14'b0000101_0000100;
		logarithm_table[4187] = 14'b0000101_0000100;
		logarithm_table[4188] = 14'b0000101_0000100;
		logarithm_table[4189] = 14'b0000101_0000100;
		logarithm_table[4190] = 14'b0000101_0000100;
		logarithm_table[4191] = 14'b0000101_0000100;
		logarithm_table[4192] = 14'b0000101_0000100;
		logarithm_table[4193] = 14'b0000101_0000100;
		logarithm_table[4194] = 14'b0000101_0000100;
		logarithm_table[4195] = 14'b0000101_0000100;
		logarithm_table[4196] = 14'b0000101_0000100;
		logarithm_table[4197] = 14'b0000101_0000100;
		logarithm_table[4198] = 14'b0000101_0000101;
		logarithm_table[4199] = 14'b0000101_0000101;
		logarithm_table[4200] = 14'b0000101_0000101;
		logarithm_table[4201] = 14'b0000101_0000101;
		logarithm_table[4202] = 14'b0000101_0000101;
		logarithm_table[4203] = 14'b0000101_0000101;
		logarithm_table[4204] = 14'b0000101_0000101;
		logarithm_table[4205] = 14'b0000101_0000101;
		logarithm_table[4206] = 14'b0000101_0000101;
		logarithm_table[4207] = 14'b0000101_0000101;
		logarithm_table[4208] = 14'b0000101_0000101;
		logarithm_table[4209] = 14'b0000101_0000101;
		logarithm_table[4210] = 14'b0000101_0000101;
		logarithm_table[4211] = 14'b0000101_0000101;
		logarithm_table[4212] = 14'b0000101_0000101;
		logarithm_table[4213] = 14'b0000101_0000101;
		logarithm_table[4214] = 14'b0000101_0000101;
		logarithm_table[4215] = 14'b0000101_0000101;
		logarithm_table[4216] = 14'b0000101_0000101;
		logarithm_table[4217] = 14'b0000101_0000101;
		logarithm_table[4218] = 14'b0000101_0000101;
		logarithm_table[4219] = 14'b0000101_0000101;
		logarithm_table[4220] = 14'b0000101_0000110;
		logarithm_table[4221] = 14'b0000101_0000110;
		logarithm_table[4222] = 14'b0000101_0000110;
		logarithm_table[4223] = 14'b0000101_0000110;
		logarithm_table[4224] = 14'b0000101_0000110;
		logarithm_table[4225] = 14'b0000101_0000110;
		logarithm_table[4226] = 14'b0000101_0000110;
		logarithm_table[4227] = 14'b0000101_0000110;
		logarithm_table[4228] = 14'b0000101_0000110;
		logarithm_table[4229] = 14'b0000101_0000110;
		logarithm_table[4230] = 14'b0000101_0000110;
		logarithm_table[4231] = 14'b0000101_0000110;
		logarithm_table[4232] = 14'b0000101_0000110;
		logarithm_table[4233] = 14'b0000101_0000110;
		logarithm_table[4234] = 14'b0000101_0000110;
		logarithm_table[4235] = 14'b0000101_0000110;
		logarithm_table[4236] = 14'b0000101_0000110;
		logarithm_table[4237] = 14'b0000101_0000110;
		logarithm_table[4238] = 14'b0000101_0000110;
		logarithm_table[4239] = 14'b0000101_0000110;
		logarithm_table[4240] = 14'b0000101_0000110;
		logarithm_table[4241] = 14'b0000101_0000110;
		logarithm_table[4242] = 14'b0000101_0000110;
		logarithm_table[4243] = 14'b0000101_0000111;
		logarithm_table[4244] = 14'b0000101_0000111;
		logarithm_table[4245] = 14'b0000101_0000111;
		logarithm_table[4246] = 14'b0000101_0000111;
		logarithm_table[4247] = 14'b0000101_0000111;
		logarithm_table[4248] = 14'b0000101_0000111;
		logarithm_table[4249] = 14'b0000101_0000111;
		logarithm_table[4250] = 14'b0000101_0000111;
		logarithm_table[4251] = 14'b0000101_0000111;
		logarithm_table[4252] = 14'b0000101_0000111;
		logarithm_table[4253] = 14'b0000101_0000111;
		logarithm_table[4254] = 14'b0000101_0000111;
		logarithm_table[4255] = 14'b0000101_0000111;
		logarithm_table[4256] = 14'b0000101_0000111;
		logarithm_table[4257] = 14'b0000101_0000111;
		logarithm_table[4258] = 14'b0000101_0000111;
		logarithm_table[4259] = 14'b0000101_0000111;
		logarithm_table[4260] = 14'b0000101_0000111;
		logarithm_table[4261] = 14'b0000101_0000111;
		logarithm_table[4262] = 14'b0000101_0000111;
		logarithm_table[4263] = 14'b0000101_0000111;
		logarithm_table[4264] = 14'b0000101_0000111;
		logarithm_table[4265] = 14'b0000101_0000111;
		logarithm_table[4266] = 14'b0000101_0001000;
		logarithm_table[4267] = 14'b0000101_0001000;
		logarithm_table[4268] = 14'b0000101_0001000;
		logarithm_table[4269] = 14'b0000101_0001000;
		logarithm_table[4270] = 14'b0000101_0001000;
		logarithm_table[4271] = 14'b0000101_0001000;
		logarithm_table[4272] = 14'b0000101_0001000;
		logarithm_table[4273] = 14'b0000101_0001000;
		logarithm_table[4274] = 14'b0000101_0001000;
		logarithm_table[4275] = 14'b0000101_0001000;
		logarithm_table[4276] = 14'b0000101_0001000;
		logarithm_table[4277] = 14'b0000101_0001000;
		logarithm_table[4278] = 14'b0000101_0001000;
		logarithm_table[4279] = 14'b0000101_0001000;
		logarithm_table[4280] = 14'b0000101_0001000;
		logarithm_table[4281] = 14'b0000101_0001000;
		logarithm_table[4282] = 14'b0000101_0001000;
		logarithm_table[4283] = 14'b0000101_0001000;
		logarithm_table[4284] = 14'b0000101_0001000;
		logarithm_table[4285] = 14'b0000101_0001000;
		logarithm_table[4286] = 14'b0000101_0001000;
		logarithm_table[4287] = 14'b0000101_0001000;
		logarithm_table[4288] = 14'b0000101_0001000;
		logarithm_table[4289] = 14'b0000101_0001001;
		logarithm_table[4290] = 14'b0000101_0001001;
		logarithm_table[4291] = 14'b0000101_0001001;
		logarithm_table[4292] = 14'b0000101_0001001;
		logarithm_table[4293] = 14'b0000101_0001001;
		logarithm_table[4294] = 14'b0000101_0001001;
		logarithm_table[4295] = 14'b0000101_0001001;
		logarithm_table[4296] = 14'b0000101_0001001;
		logarithm_table[4297] = 14'b0000101_0001001;
		logarithm_table[4298] = 14'b0000101_0001001;
		logarithm_table[4299] = 14'b0000101_0001001;
		logarithm_table[4300] = 14'b0000101_0001001;
		logarithm_table[4301] = 14'b0000101_0001001;
		logarithm_table[4302] = 14'b0000101_0001001;
		logarithm_table[4303] = 14'b0000101_0001001;
		logarithm_table[4304] = 14'b0000101_0001001;
		logarithm_table[4305] = 14'b0000101_0001001;
		logarithm_table[4306] = 14'b0000101_0001001;
		logarithm_table[4307] = 14'b0000101_0001001;
		logarithm_table[4308] = 14'b0000101_0001001;
		logarithm_table[4309] = 14'b0000101_0001001;
		logarithm_table[4310] = 14'b0000101_0001001;
		logarithm_table[4311] = 14'b0000101_0001001;
		logarithm_table[4312] = 14'b0000101_0001001;
		logarithm_table[4313] = 14'b0000101_0001010;
		logarithm_table[4314] = 14'b0000101_0001010;
		logarithm_table[4315] = 14'b0000101_0001010;
		logarithm_table[4316] = 14'b0000101_0001010;
		logarithm_table[4317] = 14'b0000101_0001010;
		logarithm_table[4318] = 14'b0000101_0001010;
		logarithm_table[4319] = 14'b0000101_0001010;
		logarithm_table[4320] = 14'b0000101_0001010;
		logarithm_table[4321] = 14'b0000101_0001010;
		logarithm_table[4322] = 14'b0000101_0001010;
		logarithm_table[4323] = 14'b0000101_0001010;
		logarithm_table[4324] = 14'b0000101_0001010;
		logarithm_table[4325] = 14'b0000101_0001010;
		logarithm_table[4326] = 14'b0000101_0001010;
		logarithm_table[4327] = 14'b0000101_0001010;
		logarithm_table[4328] = 14'b0000101_0001010;
		logarithm_table[4329] = 14'b0000101_0001010;
		logarithm_table[4330] = 14'b0000101_0001010;
		logarithm_table[4331] = 14'b0000101_0001010;
		logarithm_table[4332] = 14'b0000101_0001010;
		logarithm_table[4333] = 14'b0000101_0001010;
		logarithm_table[4334] = 14'b0000101_0001010;
		logarithm_table[4335] = 14'b0000101_0001010;
		logarithm_table[4336] = 14'b0000101_0001011;
		logarithm_table[4337] = 14'b0000101_0001011;
		logarithm_table[4338] = 14'b0000101_0001011;
		logarithm_table[4339] = 14'b0000101_0001011;
		logarithm_table[4340] = 14'b0000101_0001011;
		logarithm_table[4341] = 14'b0000101_0001011;
		logarithm_table[4342] = 14'b0000101_0001011;
		logarithm_table[4343] = 14'b0000101_0001011;
		logarithm_table[4344] = 14'b0000101_0001011;
		logarithm_table[4345] = 14'b0000101_0001011;
		logarithm_table[4346] = 14'b0000101_0001011;
		logarithm_table[4347] = 14'b0000101_0001011;
		logarithm_table[4348] = 14'b0000101_0001011;
		logarithm_table[4349] = 14'b0000101_0001011;
		logarithm_table[4350] = 14'b0000101_0001011;
		logarithm_table[4351] = 14'b0000101_0001011;
		logarithm_table[4352] = 14'b0000101_0001011;
		logarithm_table[4353] = 14'b0000101_0001011;
		logarithm_table[4354] = 14'b0000101_0001011;
		logarithm_table[4355] = 14'b0000101_0001011;
		logarithm_table[4356] = 14'b0000101_0001011;
		logarithm_table[4357] = 14'b0000101_0001011;
		logarithm_table[4358] = 14'b0000101_0001011;
		logarithm_table[4359] = 14'b0000101_0001011;
		logarithm_table[4360] = 14'b0000101_0001100;
		logarithm_table[4361] = 14'b0000101_0001100;
		logarithm_table[4362] = 14'b0000101_0001100;
		logarithm_table[4363] = 14'b0000101_0001100;
		logarithm_table[4364] = 14'b0000101_0001100;
		logarithm_table[4365] = 14'b0000101_0001100;
		logarithm_table[4366] = 14'b0000101_0001100;
		logarithm_table[4367] = 14'b0000101_0001100;
		logarithm_table[4368] = 14'b0000101_0001100;
		logarithm_table[4369] = 14'b0000101_0001100;
		logarithm_table[4370] = 14'b0000101_0001100;
		logarithm_table[4371] = 14'b0000101_0001100;
		logarithm_table[4372] = 14'b0000101_0001100;
		logarithm_table[4373] = 14'b0000101_0001100;
		logarithm_table[4374] = 14'b0000101_0001100;
		logarithm_table[4375] = 14'b0000101_0001100;
		logarithm_table[4376] = 14'b0000101_0001100;
		logarithm_table[4377] = 14'b0000101_0001100;
		logarithm_table[4378] = 14'b0000101_0001100;
		logarithm_table[4379] = 14'b0000101_0001100;
		logarithm_table[4380] = 14'b0000101_0001100;
		logarithm_table[4381] = 14'b0000101_0001100;
		logarithm_table[4382] = 14'b0000101_0001100;
		logarithm_table[4383] = 14'b0000101_0001101;
		logarithm_table[4384] = 14'b0000101_0001101;
		logarithm_table[4385] = 14'b0000101_0001101;
		logarithm_table[4386] = 14'b0000101_0001101;
		logarithm_table[4387] = 14'b0000101_0001101;
		logarithm_table[4388] = 14'b0000101_0001101;
		logarithm_table[4389] = 14'b0000101_0001101;
		logarithm_table[4390] = 14'b0000101_0001101;
		logarithm_table[4391] = 14'b0000101_0001101;
		logarithm_table[4392] = 14'b0000101_0001101;
		logarithm_table[4393] = 14'b0000101_0001101;
		logarithm_table[4394] = 14'b0000101_0001101;
		logarithm_table[4395] = 14'b0000101_0001101;
		logarithm_table[4396] = 14'b0000101_0001101;
		logarithm_table[4397] = 14'b0000101_0001101;
		logarithm_table[4398] = 14'b0000101_0001101;
		logarithm_table[4399] = 14'b0000101_0001101;
		logarithm_table[4400] = 14'b0000101_0001101;
		logarithm_table[4401] = 14'b0000101_0001101;
		logarithm_table[4402] = 14'b0000101_0001101;
		logarithm_table[4403] = 14'b0000101_0001101;
		logarithm_table[4404] = 14'b0000101_0001101;
		logarithm_table[4405] = 14'b0000101_0001101;
		logarithm_table[4406] = 14'b0000101_0001101;
		logarithm_table[4407] = 14'b0000101_0001110;
		logarithm_table[4408] = 14'b0000101_0001110;
		logarithm_table[4409] = 14'b0000101_0001110;
		logarithm_table[4410] = 14'b0000101_0001110;
		logarithm_table[4411] = 14'b0000101_0001110;
		logarithm_table[4412] = 14'b0000101_0001110;
		logarithm_table[4413] = 14'b0000101_0001110;
		logarithm_table[4414] = 14'b0000101_0001110;
		logarithm_table[4415] = 14'b0000101_0001110;
		logarithm_table[4416] = 14'b0000101_0001110;
		logarithm_table[4417] = 14'b0000101_0001110;
		logarithm_table[4418] = 14'b0000101_0001110;
		logarithm_table[4419] = 14'b0000101_0001110;
		logarithm_table[4420] = 14'b0000101_0001110;
		logarithm_table[4421] = 14'b0000101_0001110;
		logarithm_table[4422] = 14'b0000101_0001110;
		logarithm_table[4423] = 14'b0000101_0001110;
		logarithm_table[4424] = 14'b0000101_0001110;
		logarithm_table[4425] = 14'b0000101_0001110;
		logarithm_table[4426] = 14'b0000101_0001110;
		logarithm_table[4427] = 14'b0000101_0001110;
		logarithm_table[4428] = 14'b0000101_0001110;
		logarithm_table[4429] = 14'b0000101_0001110;
		logarithm_table[4430] = 14'b0000101_0001110;
		logarithm_table[4431] = 14'b0000101_0001111;
		logarithm_table[4432] = 14'b0000101_0001111;
		logarithm_table[4433] = 14'b0000101_0001111;
		logarithm_table[4434] = 14'b0000101_0001111;
		logarithm_table[4435] = 14'b0000101_0001111;
		logarithm_table[4436] = 14'b0000101_0001111;
		logarithm_table[4437] = 14'b0000101_0001111;
		logarithm_table[4438] = 14'b0000101_0001111;
		logarithm_table[4439] = 14'b0000101_0001111;
		logarithm_table[4440] = 14'b0000101_0001111;
		logarithm_table[4441] = 14'b0000101_0001111;
		logarithm_table[4442] = 14'b0000101_0001111;
		logarithm_table[4443] = 14'b0000101_0001111;
		logarithm_table[4444] = 14'b0000101_0001111;
		logarithm_table[4445] = 14'b0000101_0001111;
		logarithm_table[4446] = 14'b0000101_0001111;
		logarithm_table[4447] = 14'b0000101_0001111;
		logarithm_table[4448] = 14'b0000101_0001111;
		logarithm_table[4449] = 14'b0000101_0001111;
		logarithm_table[4450] = 14'b0000101_0001111;
		logarithm_table[4451] = 14'b0000101_0001111;
		logarithm_table[4452] = 14'b0000101_0001111;
		logarithm_table[4453] = 14'b0000101_0001111;
		logarithm_table[4454] = 14'b0000101_0001111;
		logarithm_table[4455] = 14'b0000101_0010000;
		logarithm_table[4456] = 14'b0000101_0010000;
		logarithm_table[4457] = 14'b0000101_0010000;
		logarithm_table[4458] = 14'b0000101_0010000;
		logarithm_table[4459] = 14'b0000101_0010000;
		logarithm_table[4460] = 14'b0000101_0010000;
		logarithm_table[4461] = 14'b0000101_0010000;
		logarithm_table[4462] = 14'b0000101_0010000;
		logarithm_table[4463] = 14'b0000101_0010000;
		logarithm_table[4464] = 14'b0000101_0010000;
		logarithm_table[4465] = 14'b0000101_0010000;
		logarithm_table[4466] = 14'b0000101_0010000;
		logarithm_table[4467] = 14'b0000101_0010000;
		logarithm_table[4468] = 14'b0000101_0010000;
		logarithm_table[4469] = 14'b0000101_0010000;
		logarithm_table[4470] = 14'b0000101_0010000;
		logarithm_table[4471] = 14'b0000101_0010000;
		logarithm_table[4472] = 14'b0000101_0010000;
		logarithm_table[4473] = 14'b0000101_0010000;
		logarithm_table[4474] = 14'b0000101_0010000;
		logarithm_table[4475] = 14'b0000101_0010000;
		logarithm_table[4476] = 14'b0000101_0010000;
		logarithm_table[4477] = 14'b0000101_0010000;
		logarithm_table[4478] = 14'b0000101_0010000;
		logarithm_table[4479] = 14'b0000101_0010001;
		logarithm_table[4480] = 14'b0000101_0010001;
		logarithm_table[4481] = 14'b0000101_0010001;
		logarithm_table[4482] = 14'b0000101_0010001;
		logarithm_table[4483] = 14'b0000101_0010001;
		logarithm_table[4484] = 14'b0000101_0010001;
		logarithm_table[4485] = 14'b0000101_0010001;
		logarithm_table[4486] = 14'b0000101_0010001;
		logarithm_table[4487] = 14'b0000101_0010001;
		logarithm_table[4488] = 14'b0000101_0010001;
		logarithm_table[4489] = 14'b0000101_0010001;
		logarithm_table[4490] = 14'b0000101_0010001;
		logarithm_table[4491] = 14'b0000101_0010001;
		logarithm_table[4492] = 14'b0000101_0010001;
		logarithm_table[4493] = 14'b0000101_0010001;
		logarithm_table[4494] = 14'b0000101_0010001;
		logarithm_table[4495] = 14'b0000101_0010001;
		logarithm_table[4496] = 14'b0000101_0010001;
		logarithm_table[4497] = 14'b0000101_0010001;
		logarithm_table[4498] = 14'b0000101_0010001;
		logarithm_table[4499] = 14'b0000101_0010001;
		logarithm_table[4500] = 14'b0000101_0010001;
		logarithm_table[4501] = 14'b0000101_0010001;
		logarithm_table[4502] = 14'b0000101_0010001;
		logarithm_table[4503] = 14'b0000101_0010001;
		logarithm_table[4504] = 14'b0000101_0010010;
		logarithm_table[4505] = 14'b0000101_0010010;
		logarithm_table[4506] = 14'b0000101_0010010;
		logarithm_table[4507] = 14'b0000101_0010010;
		logarithm_table[4508] = 14'b0000101_0010010;
		logarithm_table[4509] = 14'b0000101_0010010;
		logarithm_table[4510] = 14'b0000101_0010010;
		logarithm_table[4511] = 14'b0000101_0010010;
		logarithm_table[4512] = 14'b0000101_0010010;
		logarithm_table[4513] = 14'b0000101_0010010;
		logarithm_table[4514] = 14'b0000101_0010010;
		logarithm_table[4515] = 14'b0000101_0010010;
		logarithm_table[4516] = 14'b0000101_0010010;
		logarithm_table[4517] = 14'b0000101_0010010;
		logarithm_table[4518] = 14'b0000101_0010010;
		logarithm_table[4519] = 14'b0000101_0010010;
		logarithm_table[4520] = 14'b0000101_0010010;
		logarithm_table[4521] = 14'b0000101_0010010;
		logarithm_table[4522] = 14'b0000101_0010010;
		logarithm_table[4523] = 14'b0000101_0010010;
		logarithm_table[4524] = 14'b0000101_0010010;
		logarithm_table[4525] = 14'b0000101_0010010;
		logarithm_table[4526] = 14'b0000101_0010010;
		logarithm_table[4527] = 14'b0000101_0010010;
		logarithm_table[4528] = 14'b0000101_0010011;
		logarithm_table[4529] = 14'b0000101_0010011;
		logarithm_table[4530] = 14'b0000101_0010011;
		logarithm_table[4531] = 14'b0000101_0010011;
		logarithm_table[4532] = 14'b0000101_0010011;
		logarithm_table[4533] = 14'b0000101_0010011;
		logarithm_table[4534] = 14'b0000101_0010011;
		logarithm_table[4535] = 14'b0000101_0010011;
		logarithm_table[4536] = 14'b0000101_0010011;
		logarithm_table[4537] = 14'b0000101_0010011;
		logarithm_table[4538] = 14'b0000101_0010011;
		logarithm_table[4539] = 14'b0000101_0010011;
		logarithm_table[4540] = 14'b0000101_0010011;
		logarithm_table[4541] = 14'b0000101_0010011;
		logarithm_table[4542] = 14'b0000101_0010011;
		logarithm_table[4543] = 14'b0000101_0010011;
		logarithm_table[4544] = 14'b0000101_0010011;
		logarithm_table[4545] = 14'b0000101_0010011;
		logarithm_table[4546] = 14'b0000101_0010011;
		logarithm_table[4547] = 14'b0000101_0010011;
		logarithm_table[4548] = 14'b0000101_0010011;
		logarithm_table[4549] = 14'b0000101_0010011;
		logarithm_table[4550] = 14'b0000101_0010011;
		logarithm_table[4551] = 14'b0000101_0010011;
		logarithm_table[4552] = 14'b0000101_0010011;
		logarithm_table[4553] = 14'b0000101_0010100;
		logarithm_table[4554] = 14'b0000101_0010100;
		logarithm_table[4555] = 14'b0000101_0010100;
		logarithm_table[4556] = 14'b0000101_0010100;
		logarithm_table[4557] = 14'b0000101_0010100;
		logarithm_table[4558] = 14'b0000101_0010100;
		logarithm_table[4559] = 14'b0000101_0010100;
		logarithm_table[4560] = 14'b0000101_0010100;
		logarithm_table[4561] = 14'b0000101_0010100;
		logarithm_table[4562] = 14'b0000101_0010100;
		logarithm_table[4563] = 14'b0000101_0010100;
		logarithm_table[4564] = 14'b0000101_0010100;
		logarithm_table[4565] = 14'b0000101_0010100;
		logarithm_table[4566] = 14'b0000101_0010100;
		logarithm_table[4567] = 14'b0000101_0010100;
		logarithm_table[4568] = 14'b0000101_0010100;
		logarithm_table[4569] = 14'b0000101_0010100;
		logarithm_table[4570] = 14'b0000101_0010100;
		logarithm_table[4571] = 14'b0000101_0010100;
		logarithm_table[4572] = 14'b0000101_0010100;
		logarithm_table[4573] = 14'b0000101_0010100;
		logarithm_table[4574] = 14'b0000101_0010100;
		logarithm_table[4575] = 14'b0000101_0010100;
		logarithm_table[4576] = 14'b0000101_0010100;
		logarithm_table[4577] = 14'b0000101_0010101;
		logarithm_table[4578] = 14'b0000101_0010101;
		logarithm_table[4579] = 14'b0000101_0010101;
		logarithm_table[4580] = 14'b0000101_0010101;
		logarithm_table[4581] = 14'b0000101_0010101;
		logarithm_table[4582] = 14'b0000101_0010101;
		logarithm_table[4583] = 14'b0000101_0010101;
		logarithm_table[4584] = 14'b0000101_0010101;
		logarithm_table[4585] = 14'b0000101_0010101;
		logarithm_table[4586] = 14'b0000101_0010101;
		logarithm_table[4587] = 14'b0000101_0010101;
		logarithm_table[4588] = 14'b0000101_0010101;
		logarithm_table[4589] = 14'b0000101_0010101;
		logarithm_table[4590] = 14'b0000101_0010101;
		logarithm_table[4591] = 14'b0000101_0010101;
		logarithm_table[4592] = 14'b0000101_0010101;
		logarithm_table[4593] = 14'b0000101_0010101;
		logarithm_table[4594] = 14'b0000101_0010101;
		logarithm_table[4595] = 14'b0000101_0010101;
		logarithm_table[4596] = 14'b0000101_0010101;
		logarithm_table[4597] = 14'b0000101_0010101;
		logarithm_table[4598] = 14'b0000101_0010101;
		logarithm_table[4599] = 14'b0000101_0010101;
		logarithm_table[4600] = 14'b0000101_0010101;
		logarithm_table[4601] = 14'b0000101_0010101;
		logarithm_table[4602] = 14'b0000101_0010110;
		logarithm_table[4603] = 14'b0000101_0010110;
		logarithm_table[4604] = 14'b0000101_0010110;
		logarithm_table[4605] = 14'b0000101_0010110;
		logarithm_table[4606] = 14'b0000101_0010110;
		logarithm_table[4607] = 14'b0000101_0010110;
		logarithm_table[4608] = 14'b0000101_0010110;
		logarithm_table[4609] = 14'b0000101_0010110;
		logarithm_table[4610] = 14'b0000101_0010110;
		logarithm_table[4611] = 14'b0000101_0010110;
		logarithm_table[4612] = 14'b0000101_0010110;
		logarithm_table[4613] = 14'b0000101_0010110;
		logarithm_table[4614] = 14'b0000101_0010110;
		logarithm_table[4615] = 14'b0000101_0010110;
		logarithm_table[4616] = 14'b0000101_0010110;
		logarithm_table[4617] = 14'b0000101_0010110;
		logarithm_table[4618] = 14'b0000101_0010110;
		logarithm_table[4619] = 14'b0000101_0010110;
		logarithm_table[4620] = 14'b0000101_0010110;
		logarithm_table[4621] = 14'b0000101_0010110;
		logarithm_table[4622] = 14'b0000101_0010110;
		logarithm_table[4623] = 14'b0000101_0010110;
		logarithm_table[4624] = 14'b0000101_0010110;
		logarithm_table[4625] = 14'b0000101_0010110;
		logarithm_table[4626] = 14'b0000101_0010110;
		logarithm_table[4627] = 14'b0000101_0010111;
		logarithm_table[4628] = 14'b0000101_0010111;
		logarithm_table[4629] = 14'b0000101_0010111;
		logarithm_table[4630] = 14'b0000101_0010111;
		logarithm_table[4631] = 14'b0000101_0010111;
		logarithm_table[4632] = 14'b0000101_0010111;
		logarithm_table[4633] = 14'b0000101_0010111;
		logarithm_table[4634] = 14'b0000101_0010111;
		logarithm_table[4635] = 14'b0000101_0010111;
		logarithm_table[4636] = 14'b0000101_0010111;
		logarithm_table[4637] = 14'b0000101_0010111;
		logarithm_table[4638] = 14'b0000101_0010111;
		logarithm_table[4639] = 14'b0000101_0010111;
		logarithm_table[4640] = 14'b0000101_0010111;
		logarithm_table[4641] = 14'b0000101_0010111;
		logarithm_table[4642] = 14'b0000101_0010111;
		logarithm_table[4643] = 14'b0000101_0010111;
		logarithm_table[4644] = 14'b0000101_0010111;
		logarithm_table[4645] = 14'b0000101_0010111;
		logarithm_table[4646] = 14'b0000101_0010111;
		logarithm_table[4647] = 14'b0000101_0010111;
		logarithm_table[4648] = 14'b0000101_0010111;
		logarithm_table[4649] = 14'b0000101_0010111;
		logarithm_table[4650] = 14'b0000101_0010111;
		logarithm_table[4651] = 14'b0000101_0010111;
		logarithm_table[4652] = 14'b0000101_0011000;
		logarithm_table[4653] = 14'b0000101_0011000;
		logarithm_table[4654] = 14'b0000101_0011000;
		logarithm_table[4655] = 14'b0000101_0011000;
		logarithm_table[4656] = 14'b0000101_0011000;
		logarithm_table[4657] = 14'b0000101_0011000;
		logarithm_table[4658] = 14'b0000101_0011000;
		logarithm_table[4659] = 14'b0000101_0011000;
		logarithm_table[4660] = 14'b0000101_0011000;
		logarithm_table[4661] = 14'b0000101_0011000;
		logarithm_table[4662] = 14'b0000101_0011000;
		logarithm_table[4663] = 14'b0000101_0011000;
		logarithm_table[4664] = 14'b0000101_0011000;
		logarithm_table[4665] = 14'b0000101_0011000;
		logarithm_table[4666] = 14'b0000101_0011000;
		logarithm_table[4667] = 14'b0000101_0011000;
		logarithm_table[4668] = 14'b0000101_0011000;
		logarithm_table[4669] = 14'b0000101_0011000;
		logarithm_table[4670] = 14'b0000101_0011000;
		logarithm_table[4671] = 14'b0000101_0011000;
		logarithm_table[4672] = 14'b0000101_0011000;
		logarithm_table[4673] = 14'b0000101_0011000;
		logarithm_table[4674] = 14'b0000101_0011000;
		logarithm_table[4675] = 14'b0000101_0011000;
		logarithm_table[4676] = 14'b0000101_0011000;
		logarithm_table[4677] = 14'b0000101_0011000;
		logarithm_table[4678] = 14'b0000101_0011001;
		logarithm_table[4679] = 14'b0000101_0011001;
		logarithm_table[4680] = 14'b0000101_0011001;
		logarithm_table[4681] = 14'b0000101_0011001;
		logarithm_table[4682] = 14'b0000101_0011001;
		logarithm_table[4683] = 14'b0000101_0011001;
		logarithm_table[4684] = 14'b0000101_0011001;
		logarithm_table[4685] = 14'b0000101_0011001;
		logarithm_table[4686] = 14'b0000101_0011001;
		logarithm_table[4687] = 14'b0000101_0011001;
		logarithm_table[4688] = 14'b0000101_0011001;
		logarithm_table[4689] = 14'b0000101_0011001;
		logarithm_table[4690] = 14'b0000101_0011001;
		logarithm_table[4691] = 14'b0000101_0011001;
		logarithm_table[4692] = 14'b0000101_0011001;
		logarithm_table[4693] = 14'b0000101_0011001;
		logarithm_table[4694] = 14'b0000101_0011001;
		logarithm_table[4695] = 14'b0000101_0011001;
		logarithm_table[4696] = 14'b0000101_0011001;
		logarithm_table[4697] = 14'b0000101_0011001;
		logarithm_table[4698] = 14'b0000101_0011001;
		logarithm_table[4699] = 14'b0000101_0011001;
		logarithm_table[4700] = 14'b0000101_0011001;
		logarithm_table[4701] = 14'b0000101_0011001;
		logarithm_table[4702] = 14'b0000101_0011001;
		logarithm_table[4703] = 14'b0000101_0011010;
		logarithm_table[4704] = 14'b0000101_0011010;
		logarithm_table[4705] = 14'b0000101_0011010;
		logarithm_table[4706] = 14'b0000101_0011010;
		logarithm_table[4707] = 14'b0000101_0011010;
		logarithm_table[4708] = 14'b0000101_0011010;
		logarithm_table[4709] = 14'b0000101_0011010;
		logarithm_table[4710] = 14'b0000101_0011010;
		logarithm_table[4711] = 14'b0000101_0011010;
		logarithm_table[4712] = 14'b0000101_0011010;
		logarithm_table[4713] = 14'b0000101_0011010;
		logarithm_table[4714] = 14'b0000101_0011010;
		logarithm_table[4715] = 14'b0000101_0011010;
		logarithm_table[4716] = 14'b0000101_0011010;
		logarithm_table[4717] = 14'b0000101_0011010;
		logarithm_table[4718] = 14'b0000101_0011010;
		logarithm_table[4719] = 14'b0000101_0011010;
		logarithm_table[4720] = 14'b0000101_0011010;
		logarithm_table[4721] = 14'b0000101_0011010;
		logarithm_table[4722] = 14'b0000101_0011010;
		logarithm_table[4723] = 14'b0000101_0011010;
		logarithm_table[4724] = 14'b0000101_0011010;
		logarithm_table[4725] = 14'b0000101_0011010;
		logarithm_table[4726] = 14'b0000101_0011010;
		logarithm_table[4727] = 14'b0000101_0011010;
		logarithm_table[4728] = 14'b0000101_0011010;
		logarithm_table[4729] = 14'b0000101_0011011;
		logarithm_table[4730] = 14'b0000101_0011011;
		logarithm_table[4731] = 14'b0000101_0011011;
		logarithm_table[4732] = 14'b0000101_0011011;
		logarithm_table[4733] = 14'b0000101_0011011;
		logarithm_table[4734] = 14'b0000101_0011011;
		logarithm_table[4735] = 14'b0000101_0011011;
		logarithm_table[4736] = 14'b0000101_0011011;
		logarithm_table[4737] = 14'b0000101_0011011;
		logarithm_table[4738] = 14'b0000101_0011011;
		logarithm_table[4739] = 14'b0000101_0011011;
		logarithm_table[4740] = 14'b0000101_0011011;
		logarithm_table[4741] = 14'b0000101_0011011;
		logarithm_table[4742] = 14'b0000101_0011011;
		logarithm_table[4743] = 14'b0000101_0011011;
		logarithm_table[4744] = 14'b0000101_0011011;
		logarithm_table[4745] = 14'b0000101_0011011;
		logarithm_table[4746] = 14'b0000101_0011011;
		logarithm_table[4747] = 14'b0000101_0011011;
		logarithm_table[4748] = 14'b0000101_0011011;
		logarithm_table[4749] = 14'b0000101_0011011;
		logarithm_table[4750] = 14'b0000101_0011011;
		logarithm_table[4751] = 14'b0000101_0011011;
		logarithm_table[4752] = 14'b0000101_0011011;
		logarithm_table[4753] = 14'b0000101_0011011;
		logarithm_table[4754] = 14'b0000101_0011100;
		logarithm_table[4755] = 14'b0000101_0011100;
		logarithm_table[4756] = 14'b0000101_0011100;
		logarithm_table[4757] = 14'b0000101_0011100;
		logarithm_table[4758] = 14'b0000101_0011100;
		logarithm_table[4759] = 14'b0000101_0011100;
		logarithm_table[4760] = 14'b0000101_0011100;
		logarithm_table[4761] = 14'b0000101_0011100;
		logarithm_table[4762] = 14'b0000101_0011100;
		logarithm_table[4763] = 14'b0000101_0011100;
		logarithm_table[4764] = 14'b0000101_0011100;
		logarithm_table[4765] = 14'b0000101_0011100;
		logarithm_table[4766] = 14'b0000101_0011100;
		logarithm_table[4767] = 14'b0000101_0011100;
		logarithm_table[4768] = 14'b0000101_0011100;
		logarithm_table[4769] = 14'b0000101_0011100;
		logarithm_table[4770] = 14'b0000101_0011100;
		logarithm_table[4771] = 14'b0000101_0011100;
		logarithm_table[4772] = 14'b0000101_0011100;
		logarithm_table[4773] = 14'b0000101_0011100;
		logarithm_table[4774] = 14'b0000101_0011100;
		logarithm_table[4775] = 14'b0000101_0011100;
		logarithm_table[4776] = 14'b0000101_0011100;
		logarithm_table[4777] = 14'b0000101_0011100;
		logarithm_table[4778] = 14'b0000101_0011100;
		logarithm_table[4779] = 14'b0000101_0011100;
		logarithm_table[4780] = 14'b0000101_0011101;
		logarithm_table[4781] = 14'b0000101_0011101;
		logarithm_table[4782] = 14'b0000101_0011101;
		logarithm_table[4783] = 14'b0000101_0011101;
		logarithm_table[4784] = 14'b0000101_0011101;
		logarithm_table[4785] = 14'b0000101_0011101;
		logarithm_table[4786] = 14'b0000101_0011101;
		logarithm_table[4787] = 14'b0000101_0011101;
		logarithm_table[4788] = 14'b0000101_0011101;
		logarithm_table[4789] = 14'b0000101_0011101;
		logarithm_table[4790] = 14'b0000101_0011101;
		logarithm_table[4791] = 14'b0000101_0011101;
		logarithm_table[4792] = 14'b0000101_0011101;
		logarithm_table[4793] = 14'b0000101_0011101;
		logarithm_table[4794] = 14'b0000101_0011101;
		logarithm_table[4795] = 14'b0000101_0011101;
		logarithm_table[4796] = 14'b0000101_0011101;
		logarithm_table[4797] = 14'b0000101_0011101;
		logarithm_table[4798] = 14'b0000101_0011101;
		logarithm_table[4799] = 14'b0000101_0011101;
		logarithm_table[4800] = 14'b0000101_0011101;
		logarithm_table[4801] = 14'b0000101_0011101;
		logarithm_table[4802] = 14'b0000101_0011101;
		logarithm_table[4803] = 14'b0000101_0011101;
		logarithm_table[4804] = 14'b0000101_0011101;
		logarithm_table[4805] = 14'b0000101_0011101;
		logarithm_table[4806] = 14'b0000101_0011110;
		logarithm_table[4807] = 14'b0000101_0011110;
		logarithm_table[4808] = 14'b0000101_0011110;
		logarithm_table[4809] = 14'b0000101_0011110;
		logarithm_table[4810] = 14'b0000101_0011110;
		logarithm_table[4811] = 14'b0000101_0011110;
		logarithm_table[4812] = 14'b0000101_0011110;
		logarithm_table[4813] = 14'b0000101_0011110;
		logarithm_table[4814] = 14'b0000101_0011110;
		logarithm_table[4815] = 14'b0000101_0011110;
		logarithm_table[4816] = 14'b0000101_0011110;
		logarithm_table[4817] = 14'b0000101_0011110;
		logarithm_table[4818] = 14'b0000101_0011110;
		logarithm_table[4819] = 14'b0000101_0011110;
		logarithm_table[4820] = 14'b0000101_0011110;
		logarithm_table[4821] = 14'b0000101_0011110;
		logarithm_table[4822] = 14'b0000101_0011110;
		logarithm_table[4823] = 14'b0000101_0011110;
		logarithm_table[4824] = 14'b0000101_0011110;
		logarithm_table[4825] = 14'b0000101_0011110;
		logarithm_table[4826] = 14'b0000101_0011110;
		logarithm_table[4827] = 14'b0000101_0011110;
		logarithm_table[4828] = 14'b0000101_0011110;
		logarithm_table[4829] = 14'b0000101_0011110;
		logarithm_table[4830] = 14'b0000101_0011110;
		logarithm_table[4831] = 14'b0000101_0011110;
		logarithm_table[4832] = 14'b0000101_0011111;
		logarithm_table[4833] = 14'b0000101_0011111;
		logarithm_table[4834] = 14'b0000101_0011111;
		logarithm_table[4835] = 14'b0000101_0011111;
		logarithm_table[4836] = 14'b0000101_0011111;
		logarithm_table[4837] = 14'b0000101_0011111;
		logarithm_table[4838] = 14'b0000101_0011111;
		logarithm_table[4839] = 14'b0000101_0011111;
		logarithm_table[4840] = 14'b0000101_0011111;
		logarithm_table[4841] = 14'b0000101_0011111;
		logarithm_table[4842] = 14'b0000101_0011111;
		logarithm_table[4843] = 14'b0000101_0011111;
		logarithm_table[4844] = 14'b0000101_0011111;
		logarithm_table[4845] = 14'b0000101_0011111;
		logarithm_table[4846] = 14'b0000101_0011111;
		logarithm_table[4847] = 14'b0000101_0011111;
		logarithm_table[4848] = 14'b0000101_0011111;
		logarithm_table[4849] = 14'b0000101_0011111;
		logarithm_table[4850] = 14'b0000101_0011111;
		logarithm_table[4851] = 14'b0000101_0011111;
		logarithm_table[4852] = 14'b0000101_0011111;
		logarithm_table[4853] = 14'b0000101_0011111;
		logarithm_table[4854] = 14'b0000101_0011111;
		logarithm_table[4855] = 14'b0000101_0011111;
		logarithm_table[4856] = 14'b0000101_0011111;
		logarithm_table[4857] = 14'b0000101_0011111;
		logarithm_table[4858] = 14'b0000101_0100000;
		logarithm_table[4859] = 14'b0000101_0100000;
		logarithm_table[4860] = 14'b0000101_0100000;
		logarithm_table[4861] = 14'b0000101_0100000;
		logarithm_table[4862] = 14'b0000101_0100000;
		logarithm_table[4863] = 14'b0000101_0100000;
		logarithm_table[4864] = 14'b0000101_0100000;
		logarithm_table[4865] = 14'b0000101_0100000;
		logarithm_table[4866] = 14'b0000101_0100000;
		logarithm_table[4867] = 14'b0000101_0100000;
		logarithm_table[4868] = 14'b0000101_0100000;
		logarithm_table[4869] = 14'b0000101_0100000;
		logarithm_table[4870] = 14'b0000101_0100000;
		logarithm_table[4871] = 14'b0000101_0100000;
		logarithm_table[4872] = 14'b0000101_0100000;
		logarithm_table[4873] = 14'b0000101_0100000;
		logarithm_table[4874] = 14'b0000101_0100000;
		logarithm_table[4875] = 14'b0000101_0100000;
		logarithm_table[4876] = 14'b0000101_0100000;
		logarithm_table[4877] = 14'b0000101_0100000;
		logarithm_table[4878] = 14'b0000101_0100000;
		logarithm_table[4879] = 14'b0000101_0100000;
		logarithm_table[4880] = 14'b0000101_0100000;
		logarithm_table[4881] = 14'b0000101_0100000;
		logarithm_table[4882] = 14'b0000101_0100000;
		logarithm_table[4883] = 14'b0000101_0100000;
		logarithm_table[4884] = 14'b0000101_0100000;
		logarithm_table[4885] = 14'b0000101_0100001;
		logarithm_table[4886] = 14'b0000101_0100001;
		logarithm_table[4887] = 14'b0000101_0100001;
		logarithm_table[4888] = 14'b0000101_0100001;
		logarithm_table[4889] = 14'b0000101_0100001;
		logarithm_table[4890] = 14'b0000101_0100001;
		logarithm_table[4891] = 14'b0000101_0100001;
		logarithm_table[4892] = 14'b0000101_0100001;
		logarithm_table[4893] = 14'b0000101_0100001;
		logarithm_table[4894] = 14'b0000101_0100001;
		logarithm_table[4895] = 14'b0000101_0100001;
		logarithm_table[4896] = 14'b0000101_0100001;
		logarithm_table[4897] = 14'b0000101_0100001;
		logarithm_table[4898] = 14'b0000101_0100001;
		logarithm_table[4899] = 14'b0000101_0100001;
		logarithm_table[4900] = 14'b0000101_0100001;
		logarithm_table[4901] = 14'b0000101_0100001;
		logarithm_table[4902] = 14'b0000101_0100001;
		logarithm_table[4903] = 14'b0000101_0100001;
		logarithm_table[4904] = 14'b0000101_0100001;
		logarithm_table[4905] = 14'b0000101_0100001;
		logarithm_table[4906] = 14'b0000101_0100001;
		logarithm_table[4907] = 14'b0000101_0100001;
		logarithm_table[4908] = 14'b0000101_0100001;
		logarithm_table[4909] = 14'b0000101_0100001;
		logarithm_table[4910] = 14'b0000101_0100001;
		logarithm_table[4911] = 14'b0000101_0100010;
		logarithm_table[4912] = 14'b0000101_0100010;
		logarithm_table[4913] = 14'b0000101_0100010;
		logarithm_table[4914] = 14'b0000101_0100010;
		logarithm_table[4915] = 14'b0000101_0100010;
		logarithm_table[4916] = 14'b0000101_0100010;
		logarithm_table[4917] = 14'b0000101_0100010;
		logarithm_table[4918] = 14'b0000101_0100010;
		logarithm_table[4919] = 14'b0000101_0100010;
		logarithm_table[4920] = 14'b0000101_0100010;
		logarithm_table[4921] = 14'b0000101_0100010;
		logarithm_table[4922] = 14'b0000101_0100010;
		logarithm_table[4923] = 14'b0000101_0100010;
		logarithm_table[4924] = 14'b0000101_0100010;
		logarithm_table[4925] = 14'b0000101_0100010;
		logarithm_table[4926] = 14'b0000101_0100010;
		logarithm_table[4927] = 14'b0000101_0100010;
		logarithm_table[4928] = 14'b0000101_0100010;
		logarithm_table[4929] = 14'b0000101_0100010;
		logarithm_table[4930] = 14'b0000101_0100010;
		logarithm_table[4931] = 14'b0000101_0100010;
		logarithm_table[4932] = 14'b0000101_0100010;
		logarithm_table[4933] = 14'b0000101_0100010;
		logarithm_table[4934] = 14'b0000101_0100010;
		logarithm_table[4935] = 14'b0000101_0100010;
		logarithm_table[4936] = 14'b0000101_0100010;
		logarithm_table[4937] = 14'b0000101_0100010;
		logarithm_table[4938] = 14'b0000101_0100011;
		logarithm_table[4939] = 14'b0000101_0100011;
		logarithm_table[4940] = 14'b0000101_0100011;
		logarithm_table[4941] = 14'b0000101_0100011;
		logarithm_table[4942] = 14'b0000101_0100011;
		logarithm_table[4943] = 14'b0000101_0100011;
		logarithm_table[4944] = 14'b0000101_0100011;
		logarithm_table[4945] = 14'b0000101_0100011;
		logarithm_table[4946] = 14'b0000101_0100011;
		logarithm_table[4947] = 14'b0000101_0100011;
		logarithm_table[4948] = 14'b0000101_0100011;
		logarithm_table[4949] = 14'b0000101_0100011;
		logarithm_table[4950] = 14'b0000101_0100011;
		logarithm_table[4951] = 14'b0000101_0100011;
		logarithm_table[4952] = 14'b0000101_0100011;
		logarithm_table[4953] = 14'b0000101_0100011;
		logarithm_table[4954] = 14'b0000101_0100011;
		logarithm_table[4955] = 14'b0000101_0100011;
		logarithm_table[4956] = 14'b0000101_0100011;
		logarithm_table[4957] = 14'b0000101_0100011;
		logarithm_table[4958] = 14'b0000101_0100011;
		logarithm_table[4959] = 14'b0000101_0100011;
		logarithm_table[4960] = 14'b0000101_0100011;
		logarithm_table[4961] = 14'b0000101_0100011;
		logarithm_table[4962] = 14'b0000101_0100011;
		logarithm_table[4963] = 14'b0000101_0100011;
		logarithm_table[4964] = 14'b0000101_0100011;
		logarithm_table[4965] = 14'b0000101_0100100;
		logarithm_table[4966] = 14'b0000101_0100100;
		logarithm_table[4967] = 14'b0000101_0100100;
		logarithm_table[4968] = 14'b0000101_0100100;
		logarithm_table[4969] = 14'b0000101_0100100;
		logarithm_table[4970] = 14'b0000101_0100100;
		logarithm_table[4971] = 14'b0000101_0100100;
		logarithm_table[4972] = 14'b0000101_0100100;
		logarithm_table[4973] = 14'b0000101_0100100;
		logarithm_table[4974] = 14'b0000101_0100100;
		logarithm_table[4975] = 14'b0000101_0100100;
		logarithm_table[4976] = 14'b0000101_0100100;
		logarithm_table[4977] = 14'b0000101_0100100;
		logarithm_table[4978] = 14'b0000101_0100100;
		logarithm_table[4979] = 14'b0000101_0100100;
		logarithm_table[4980] = 14'b0000101_0100100;
		logarithm_table[4981] = 14'b0000101_0100100;
		logarithm_table[4982] = 14'b0000101_0100100;
		logarithm_table[4983] = 14'b0000101_0100100;
		logarithm_table[4984] = 14'b0000101_0100100;
		logarithm_table[4985] = 14'b0000101_0100100;
		logarithm_table[4986] = 14'b0000101_0100100;
		logarithm_table[4987] = 14'b0000101_0100100;
		logarithm_table[4988] = 14'b0000101_0100100;
		logarithm_table[4989] = 14'b0000101_0100100;
		logarithm_table[4990] = 14'b0000101_0100100;
		logarithm_table[4991] = 14'b0000101_0100100;
		logarithm_table[4992] = 14'b0000101_0100101;
		logarithm_table[4993] = 14'b0000101_0100101;
		logarithm_table[4994] = 14'b0000101_0100101;
		logarithm_table[4995] = 14'b0000101_0100101;
		logarithm_table[4996] = 14'b0000101_0100101;
		logarithm_table[4997] = 14'b0000101_0100101;
		logarithm_table[4998] = 14'b0000101_0100101;
		logarithm_table[4999] = 14'b0000101_0100101;
		logarithm_table[5000] = 14'b0000101_0100101;
		logarithm_table[5001] = 14'b0000101_0100101;
		logarithm_table[5002] = 14'b0000101_0100101;
		logarithm_table[5003] = 14'b0000101_0100101;
		logarithm_table[5004] = 14'b0000101_0100101;
		logarithm_table[5005] = 14'b0000101_0100101;
		logarithm_table[5006] = 14'b0000101_0100101;
		logarithm_table[5007] = 14'b0000101_0100101;
		logarithm_table[5008] = 14'b0000101_0100101;
		logarithm_table[5009] = 14'b0000101_0100101;
		logarithm_table[5010] = 14'b0000101_0100101;
		logarithm_table[5011] = 14'b0000101_0100101;
		logarithm_table[5012] = 14'b0000101_0100101;
		logarithm_table[5013] = 14'b0000101_0100101;
		logarithm_table[5014] = 14'b0000101_0100101;
		logarithm_table[5015] = 14'b0000101_0100101;
		logarithm_table[5016] = 14'b0000101_0100101;
		logarithm_table[5017] = 14'b0000101_0100101;
		logarithm_table[5018] = 14'b0000101_0100101;
		logarithm_table[5019] = 14'b0000101_0100110;
		logarithm_table[5020] = 14'b0000101_0100110;
		logarithm_table[5021] = 14'b0000101_0100110;
		logarithm_table[5022] = 14'b0000101_0100110;
		logarithm_table[5023] = 14'b0000101_0100110;
		logarithm_table[5024] = 14'b0000101_0100110;
		logarithm_table[5025] = 14'b0000101_0100110;
		logarithm_table[5026] = 14'b0000101_0100110;
		logarithm_table[5027] = 14'b0000101_0100110;
		logarithm_table[5028] = 14'b0000101_0100110;
		logarithm_table[5029] = 14'b0000101_0100110;
		logarithm_table[5030] = 14'b0000101_0100110;
		logarithm_table[5031] = 14'b0000101_0100110;
		logarithm_table[5032] = 14'b0000101_0100110;
		logarithm_table[5033] = 14'b0000101_0100110;
		logarithm_table[5034] = 14'b0000101_0100110;
		logarithm_table[5035] = 14'b0000101_0100110;
		logarithm_table[5036] = 14'b0000101_0100110;
		logarithm_table[5037] = 14'b0000101_0100110;
		logarithm_table[5038] = 14'b0000101_0100110;
		logarithm_table[5039] = 14'b0000101_0100110;
		logarithm_table[5040] = 14'b0000101_0100110;
		logarithm_table[5041] = 14'b0000101_0100110;
		logarithm_table[5042] = 14'b0000101_0100110;
		logarithm_table[5043] = 14'b0000101_0100110;
		logarithm_table[5044] = 14'b0000101_0100110;
		logarithm_table[5045] = 14'b0000101_0100110;
		logarithm_table[5046] = 14'b0000101_0100111;
		logarithm_table[5047] = 14'b0000101_0100111;
		logarithm_table[5048] = 14'b0000101_0100111;
		logarithm_table[5049] = 14'b0000101_0100111;
		logarithm_table[5050] = 14'b0000101_0100111;
		logarithm_table[5051] = 14'b0000101_0100111;
		logarithm_table[5052] = 14'b0000101_0100111;
		logarithm_table[5053] = 14'b0000101_0100111;
		logarithm_table[5054] = 14'b0000101_0100111;
		logarithm_table[5055] = 14'b0000101_0100111;
		logarithm_table[5056] = 14'b0000101_0100111;
		logarithm_table[5057] = 14'b0000101_0100111;
		logarithm_table[5058] = 14'b0000101_0100111;
		logarithm_table[5059] = 14'b0000101_0100111;
		logarithm_table[5060] = 14'b0000101_0100111;
		logarithm_table[5061] = 14'b0000101_0100111;
		logarithm_table[5062] = 14'b0000101_0100111;
		logarithm_table[5063] = 14'b0000101_0100111;
		logarithm_table[5064] = 14'b0000101_0100111;
		logarithm_table[5065] = 14'b0000101_0100111;
		logarithm_table[5066] = 14'b0000101_0100111;
		logarithm_table[5067] = 14'b0000101_0100111;
		logarithm_table[5068] = 14'b0000101_0100111;
		logarithm_table[5069] = 14'b0000101_0100111;
		logarithm_table[5070] = 14'b0000101_0100111;
		logarithm_table[5071] = 14'b0000101_0100111;
		logarithm_table[5072] = 14'b0000101_0100111;
		logarithm_table[5073] = 14'b0000101_0101000;
		logarithm_table[5074] = 14'b0000101_0101000;
		logarithm_table[5075] = 14'b0000101_0101000;
		logarithm_table[5076] = 14'b0000101_0101000;
		logarithm_table[5077] = 14'b0000101_0101000;
		logarithm_table[5078] = 14'b0000101_0101000;
		logarithm_table[5079] = 14'b0000101_0101000;
		logarithm_table[5080] = 14'b0000101_0101000;
		logarithm_table[5081] = 14'b0000101_0101000;
		logarithm_table[5082] = 14'b0000101_0101000;
		logarithm_table[5083] = 14'b0000101_0101000;
		logarithm_table[5084] = 14'b0000101_0101000;
		logarithm_table[5085] = 14'b0000101_0101000;
		logarithm_table[5086] = 14'b0000101_0101000;
		logarithm_table[5087] = 14'b0000101_0101000;
		logarithm_table[5088] = 14'b0000101_0101000;
		logarithm_table[5089] = 14'b0000101_0101000;
		logarithm_table[5090] = 14'b0000101_0101000;
		logarithm_table[5091] = 14'b0000101_0101000;
		logarithm_table[5092] = 14'b0000101_0101000;
		logarithm_table[5093] = 14'b0000101_0101000;
		logarithm_table[5094] = 14'b0000101_0101000;
		logarithm_table[5095] = 14'b0000101_0101000;
		logarithm_table[5096] = 14'b0000101_0101000;
		logarithm_table[5097] = 14'b0000101_0101000;
		logarithm_table[5098] = 14'b0000101_0101000;
		logarithm_table[5099] = 14'b0000101_0101000;
		logarithm_table[5100] = 14'b0000101_0101000;
		logarithm_table[5101] = 14'b0000101_0101001;
		logarithm_table[5102] = 14'b0000101_0101001;
		logarithm_table[5103] = 14'b0000101_0101001;
		logarithm_table[5104] = 14'b0000101_0101001;
		logarithm_table[5105] = 14'b0000101_0101001;
		logarithm_table[5106] = 14'b0000101_0101001;
		logarithm_table[5107] = 14'b0000101_0101001;
		logarithm_table[5108] = 14'b0000101_0101001;
		logarithm_table[5109] = 14'b0000101_0101001;
		logarithm_table[5110] = 14'b0000101_0101001;
		logarithm_table[5111] = 14'b0000101_0101001;
		logarithm_table[5112] = 14'b0000101_0101001;
		logarithm_table[5113] = 14'b0000101_0101001;
		logarithm_table[5114] = 14'b0000101_0101001;
		logarithm_table[5115] = 14'b0000101_0101001;
		logarithm_table[5116] = 14'b0000101_0101001;
		logarithm_table[5117] = 14'b0000101_0101001;
		logarithm_table[5118] = 14'b0000101_0101001;
		logarithm_table[5119] = 14'b0000101_0101001;
		logarithm_table[5120] = 14'b0000101_0101001;
		logarithm_table[5121] = 14'b0000101_0101001;
		logarithm_table[5122] = 14'b0000101_0101001;
		logarithm_table[5123] = 14'b0000101_0101001;
		logarithm_table[5124] = 14'b0000101_0101001;
		logarithm_table[5125] = 14'b0000101_0101001;
		logarithm_table[5126] = 14'b0000101_0101001;
		logarithm_table[5127] = 14'b0000101_0101001;
		logarithm_table[5128] = 14'b0000101_0101001;
		logarithm_table[5129] = 14'b0000101_0101010;
		logarithm_table[5130] = 14'b0000101_0101010;
		logarithm_table[5131] = 14'b0000101_0101010;
		logarithm_table[5132] = 14'b0000101_0101010;
		logarithm_table[5133] = 14'b0000101_0101010;
		logarithm_table[5134] = 14'b0000101_0101010;
		logarithm_table[5135] = 14'b0000101_0101010;
		logarithm_table[5136] = 14'b0000101_0101010;
		logarithm_table[5137] = 14'b0000101_0101010;
		logarithm_table[5138] = 14'b0000101_0101010;
		logarithm_table[5139] = 14'b0000101_0101010;
		logarithm_table[5140] = 14'b0000101_0101010;
		logarithm_table[5141] = 14'b0000101_0101010;
		logarithm_table[5142] = 14'b0000101_0101010;
		logarithm_table[5143] = 14'b0000101_0101010;
		logarithm_table[5144] = 14'b0000101_0101010;
		logarithm_table[5145] = 14'b0000101_0101010;
		logarithm_table[5146] = 14'b0000101_0101010;
		logarithm_table[5147] = 14'b0000101_0101010;
		logarithm_table[5148] = 14'b0000101_0101010;
		logarithm_table[5149] = 14'b0000101_0101010;
		logarithm_table[5150] = 14'b0000101_0101010;
		logarithm_table[5151] = 14'b0000101_0101010;
		logarithm_table[5152] = 14'b0000101_0101010;
		logarithm_table[5153] = 14'b0000101_0101010;
		logarithm_table[5154] = 14'b0000101_0101010;
		logarithm_table[5155] = 14'b0000101_0101010;
		logarithm_table[5156] = 14'b0000101_0101011;
		logarithm_table[5157] = 14'b0000101_0101011;
		logarithm_table[5158] = 14'b0000101_0101011;
		logarithm_table[5159] = 14'b0000101_0101011;
		logarithm_table[5160] = 14'b0000101_0101011;
		logarithm_table[5161] = 14'b0000101_0101011;
		logarithm_table[5162] = 14'b0000101_0101011;
		logarithm_table[5163] = 14'b0000101_0101011;
		logarithm_table[5164] = 14'b0000101_0101011;
		logarithm_table[5165] = 14'b0000101_0101011;
		logarithm_table[5166] = 14'b0000101_0101011;
		logarithm_table[5167] = 14'b0000101_0101011;
		logarithm_table[5168] = 14'b0000101_0101011;
		logarithm_table[5169] = 14'b0000101_0101011;
		logarithm_table[5170] = 14'b0000101_0101011;
		logarithm_table[5171] = 14'b0000101_0101011;
		logarithm_table[5172] = 14'b0000101_0101011;
		logarithm_table[5173] = 14'b0000101_0101011;
		logarithm_table[5174] = 14'b0000101_0101011;
		logarithm_table[5175] = 14'b0000101_0101011;
		logarithm_table[5176] = 14'b0000101_0101011;
		logarithm_table[5177] = 14'b0000101_0101011;
		logarithm_table[5178] = 14'b0000101_0101011;
		logarithm_table[5179] = 14'b0000101_0101011;
		logarithm_table[5180] = 14'b0000101_0101011;
		logarithm_table[5181] = 14'b0000101_0101011;
		logarithm_table[5182] = 14'b0000101_0101011;
		logarithm_table[5183] = 14'b0000101_0101011;
		logarithm_table[5184] = 14'b0000101_0101100;
		logarithm_table[5185] = 14'b0000101_0101100;
		logarithm_table[5186] = 14'b0000101_0101100;
		logarithm_table[5187] = 14'b0000101_0101100;
		logarithm_table[5188] = 14'b0000101_0101100;
		logarithm_table[5189] = 14'b0000101_0101100;
		logarithm_table[5190] = 14'b0000101_0101100;
		logarithm_table[5191] = 14'b0000101_0101100;
		logarithm_table[5192] = 14'b0000101_0101100;
		logarithm_table[5193] = 14'b0000101_0101100;
		logarithm_table[5194] = 14'b0000101_0101100;
		logarithm_table[5195] = 14'b0000101_0101100;
		logarithm_table[5196] = 14'b0000101_0101100;
		logarithm_table[5197] = 14'b0000101_0101100;
		logarithm_table[5198] = 14'b0000101_0101100;
		logarithm_table[5199] = 14'b0000101_0101100;
		logarithm_table[5200] = 14'b0000101_0101100;
		logarithm_table[5201] = 14'b0000101_0101100;
		logarithm_table[5202] = 14'b0000101_0101100;
		logarithm_table[5203] = 14'b0000101_0101100;
		logarithm_table[5204] = 14'b0000101_0101100;
		logarithm_table[5205] = 14'b0000101_0101100;
		logarithm_table[5206] = 14'b0000101_0101100;
		logarithm_table[5207] = 14'b0000101_0101100;
		logarithm_table[5208] = 14'b0000101_0101100;
		logarithm_table[5209] = 14'b0000101_0101100;
		logarithm_table[5210] = 14'b0000101_0101100;
		logarithm_table[5211] = 14'b0000101_0101100;
		logarithm_table[5212] = 14'b0000101_0101100;
		logarithm_table[5213] = 14'b0000101_0101101;
		logarithm_table[5214] = 14'b0000101_0101101;
		logarithm_table[5215] = 14'b0000101_0101101;
		logarithm_table[5216] = 14'b0000101_0101101;
		logarithm_table[5217] = 14'b0000101_0101101;
		logarithm_table[5218] = 14'b0000101_0101101;
		logarithm_table[5219] = 14'b0000101_0101101;
		logarithm_table[5220] = 14'b0000101_0101101;
		logarithm_table[5221] = 14'b0000101_0101101;
		logarithm_table[5222] = 14'b0000101_0101101;
		logarithm_table[5223] = 14'b0000101_0101101;
		logarithm_table[5224] = 14'b0000101_0101101;
		logarithm_table[5225] = 14'b0000101_0101101;
		logarithm_table[5226] = 14'b0000101_0101101;
		logarithm_table[5227] = 14'b0000101_0101101;
		logarithm_table[5228] = 14'b0000101_0101101;
		logarithm_table[5229] = 14'b0000101_0101101;
		logarithm_table[5230] = 14'b0000101_0101101;
		logarithm_table[5231] = 14'b0000101_0101101;
		logarithm_table[5232] = 14'b0000101_0101101;
		logarithm_table[5233] = 14'b0000101_0101101;
		logarithm_table[5234] = 14'b0000101_0101101;
		logarithm_table[5235] = 14'b0000101_0101101;
		logarithm_table[5236] = 14'b0000101_0101101;
		logarithm_table[5237] = 14'b0000101_0101101;
		logarithm_table[5238] = 14'b0000101_0101101;
		logarithm_table[5239] = 14'b0000101_0101101;
		logarithm_table[5240] = 14'b0000101_0101101;
		logarithm_table[5241] = 14'b0000101_0101110;
		logarithm_table[5242] = 14'b0000101_0101110;
		logarithm_table[5243] = 14'b0000101_0101110;
		logarithm_table[5244] = 14'b0000101_0101110;
		logarithm_table[5245] = 14'b0000101_0101110;
		logarithm_table[5246] = 14'b0000101_0101110;
		logarithm_table[5247] = 14'b0000101_0101110;
		logarithm_table[5248] = 14'b0000101_0101110;
		logarithm_table[5249] = 14'b0000101_0101110;
		logarithm_table[5250] = 14'b0000101_0101110;
		logarithm_table[5251] = 14'b0000101_0101110;
		logarithm_table[5252] = 14'b0000101_0101110;
		logarithm_table[5253] = 14'b0000101_0101110;
		logarithm_table[5254] = 14'b0000101_0101110;
		logarithm_table[5255] = 14'b0000101_0101110;
		logarithm_table[5256] = 14'b0000101_0101110;
		logarithm_table[5257] = 14'b0000101_0101110;
		logarithm_table[5258] = 14'b0000101_0101110;
		logarithm_table[5259] = 14'b0000101_0101110;
		logarithm_table[5260] = 14'b0000101_0101110;
		logarithm_table[5261] = 14'b0000101_0101110;
		logarithm_table[5262] = 14'b0000101_0101110;
		logarithm_table[5263] = 14'b0000101_0101110;
		logarithm_table[5264] = 14'b0000101_0101110;
		logarithm_table[5265] = 14'b0000101_0101110;
		logarithm_table[5266] = 14'b0000101_0101110;
		logarithm_table[5267] = 14'b0000101_0101110;
		logarithm_table[5268] = 14'b0000101_0101110;
		logarithm_table[5269] = 14'b0000101_0101111;
		logarithm_table[5270] = 14'b0000101_0101111;
		logarithm_table[5271] = 14'b0000101_0101111;
		logarithm_table[5272] = 14'b0000101_0101111;
		logarithm_table[5273] = 14'b0000101_0101111;
		logarithm_table[5274] = 14'b0000101_0101111;
		logarithm_table[5275] = 14'b0000101_0101111;
		logarithm_table[5276] = 14'b0000101_0101111;
		logarithm_table[5277] = 14'b0000101_0101111;
		logarithm_table[5278] = 14'b0000101_0101111;
		logarithm_table[5279] = 14'b0000101_0101111;
		logarithm_table[5280] = 14'b0000101_0101111;
		logarithm_table[5281] = 14'b0000101_0101111;
		logarithm_table[5282] = 14'b0000101_0101111;
		logarithm_table[5283] = 14'b0000101_0101111;
		logarithm_table[5284] = 14'b0000101_0101111;
		logarithm_table[5285] = 14'b0000101_0101111;
		logarithm_table[5286] = 14'b0000101_0101111;
		logarithm_table[5287] = 14'b0000101_0101111;
		logarithm_table[5288] = 14'b0000101_0101111;
		logarithm_table[5289] = 14'b0000101_0101111;
		logarithm_table[5290] = 14'b0000101_0101111;
		logarithm_table[5291] = 14'b0000101_0101111;
		logarithm_table[5292] = 14'b0000101_0101111;
		logarithm_table[5293] = 14'b0000101_0101111;
		logarithm_table[5294] = 14'b0000101_0101111;
		logarithm_table[5295] = 14'b0000101_0101111;
		logarithm_table[5296] = 14'b0000101_0101111;
		logarithm_table[5297] = 14'b0000101_0101111;
		logarithm_table[5298] = 14'b0000101_0110000;
		logarithm_table[5299] = 14'b0000101_0110000;
		logarithm_table[5300] = 14'b0000101_0110000;
		logarithm_table[5301] = 14'b0000101_0110000;
		logarithm_table[5302] = 14'b0000101_0110000;
		logarithm_table[5303] = 14'b0000101_0110000;
		logarithm_table[5304] = 14'b0000101_0110000;
		logarithm_table[5305] = 14'b0000101_0110000;
		logarithm_table[5306] = 14'b0000101_0110000;
		logarithm_table[5307] = 14'b0000101_0110000;
		logarithm_table[5308] = 14'b0000101_0110000;
		logarithm_table[5309] = 14'b0000101_0110000;
		logarithm_table[5310] = 14'b0000101_0110000;
		logarithm_table[5311] = 14'b0000101_0110000;
		logarithm_table[5312] = 14'b0000101_0110000;
		logarithm_table[5313] = 14'b0000101_0110000;
		logarithm_table[5314] = 14'b0000101_0110000;
		logarithm_table[5315] = 14'b0000101_0110000;
		logarithm_table[5316] = 14'b0000101_0110000;
		logarithm_table[5317] = 14'b0000101_0110000;
		logarithm_table[5318] = 14'b0000101_0110000;
		logarithm_table[5319] = 14'b0000101_0110000;
		logarithm_table[5320] = 14'b0000101_0110000;
		logarithm_table[5321] = 14'b0000101_0110000;
		logarithm_table[5322] = 14'b0000101_0110000;
		logarithm_table[5323] = 14'b0000101_0110000;
		logarithm_table[5324] = 14'b0000101_0110000;
		logarithm_table[5325] = 14'b0000101_0110000;
		logarithm_table[5326] = 14'b0000101_0110000;
		logarithm_table[5327] = 14'b0000101_0110001;
		logarithm_table[5328] = 14'b0000101_0110001;
		logarithm_table[5329] = 14'b0000101_0110001;
		logarithm_table[5330] = 14'b0000101_0110001;
		logarithm_table[5331] = 14'b0000101_0110001;
		logarithm_table[5332] = 14'b0000101_0110001;
		logarithm_table[5333] = 14'b0000101_0110001;
		logarithm_table[5334] = 14'b0000101_0110001;
		logarithm_table[5335] = 14'b0000101_0110001;
		logarithm_table[5336] = 14'b0000101_0110001;
		logarithm_table[5337] = 14'b0000101_0110001;
		logarithm_table[5338] = 14'b0000101_0110001;
		logarithm_table[5339] = 14'b0000101_0110001;
		logarithm_table[5340] = 14'b0000101_0110001;
		logarithm_table[5341] = 14'b0000101_0110001;
		logarithm_table[5342] = 14'b0000101_0110001;
		logarithm_table[5343] = 14'b0000101_0110001;
		logarithm_table[5344] = 14'b0000101_0110001;
		logarithm_table[5345] = 14'b0000101_0110001;
		logarithm_table[5346] = 14'b0000101_0110001;
		logarithm_table[5347] = 14'b0000101_0110001;
		logarithm_table[5348] = 14'b0000101_0110001;
		logarithm_table[5349] = 14'b0000101_0110001;
		logarithm_table[5350] = 14'b0000101_0110001;
		logarithm_table[5351] = 14'b0000101_0110001;
		logarithm_table[5352] = 14'b0000101_0110001;
		logarithm_table[5353] = 14'b0000101_0110001;
		logarithm_table[5354] = 14'b0000101_0110001;
		logarithm_table[5355] = 14'b0000101_0110001;
		logarithm_table[5356] = 14'b0000101_0110010;
		logarithm_table[5357] = 14'b0000101_0110010;
		logarithm_table[5358] = 14'b0000101_0110010;
		logarithm_table[5359] = 14'b0000101_0110010;
		logarithm_table[5360] = 14'b0000101_0110010;
		logarithm_table[5361] = 14'b0000101_0110010;
		logarithm_table[5362] = 14'b0000101_0110010;
		logarithm_table[5363] = 14'b0000101_0110010;
		logarithm_table[5364] = 14'b0000101_0110010;
		logarithm_table[5365] = 14'b0000101_0110010;
		logarithm_table[5366] = 14'b0000101_0110010;
		logarithm_table[5367] = 14'b0000101_0110010;
		logarithm_table[5368] = 14'b0000101_0110010;
		logarithm_table[5369] = 14'b0000101_0110010;
		logarithm_table[5370] = 14'b0000101_0110010;
		logarithm_table[5371] = 14'b0000101_0110010;
		logarithm_table[5372] = 14'b0000101_0110010;
		logarithm_table[5373] = 14'b0000101_0110010;
		logarithm_table[5374] = 14'b0000101_0110010;
		logarithm_table[5375] = 14'b0000101_0110010;
		logarithm_table[5376] = 14'b0000101_0110010;
		logarithm_table[5377] = 14'b0000101_0110010;
		logarithm_table[5378] = 14'b0000101_0110010;
		logarithm_table[5379] = 14'b0000101_0110010;
		logarithm_table[5380] = 14'b0000101_0110010;
		logarithm_table[5381] = 14'b0000101_0110010;
		logarithm_table[5382] = 14'b0000101_0110010;
		logarithm_table[5383] = 14'b0000101_0110010;
		logarithm_table[5384] = 14'b0000101_0110010;
		logarithm_table[5385] = 14'b0000101_0110011;
		logarithm_table[5386] = 14'b0000101_0110011;
		logarithm_table[5387] = 14'b0000101_0110011;
		logarithm_table[5388] = 14'b0000101_0110011;
		logarithm_table[5389] = 14'b0000101_0110011;
		logarithm_table[5390] = 14'b0000101_0110011;
		logarithm_table[5391] = 14'b0000101_0110011;
		logarithm_table[5392] = 14'b0000101_0110011;
		logarithm_table[5393] = 14'b0000101_0110011;
		logarithm_table[5394] = 14'b0000101_0110011;
		logarithm_table[5395] = 14'b0000101_0110011;
		logarithm_table[5396] = 14'b0000101_0110011;
		logarithm_table[5397] = 14'b0000101_0110011;
		logarithm_table[5398] = 14'b0000101_0110011;
		logarithm_table[5399] = 14'b0000101_0110011;
		logarithm_table[5400] = 14'b0000101_0110011;
		logarithm_table[5401] = 14'b0000101_0110011;
		logarithm_table[5402] = 14'b0000101_0110011;
		logarithm_table[5403] = 14'b0000101_0110011;
		logarithm_table[5404] = 14'b0000101_0110011;
		logarithm_table[5405] = 14'b0000101_0110011;
		logarithm_table[5406] = 14'b0000101_0110011;
		logarithm_table[5407] = 14'b0000101_0110011;
		logarithm_table[5408] = 14'b0000101_0110011;
		logarithm_table[5409] = 14'b0000101_0110011;
		logarithm_table[5410] = 14'b0000101_0110011;
		logarithm_table[5411] = 14'b0000101_0110011;
		logarithm_table[5412] = 14'b0000101_0110011;
		logarithm_table[5413] = 14'b0000101_0110011;
		logarithm_table[5414] = 14'b0000101_0110100;
		logarithm_table[5415] = 14'b0000101_0110100;
		logarithm_table[5416] = 14'b0000101_0110100;
		logarithm_table[5417] = 14'b0000101_0110100;
		logarithm_table[5418] = 14'b0000101_0110100;
		logarithm_table[5419] = 14'b0000101_0110100;
		logarithm_table[5420] = 14'b0000101_0110100;
		logarithm_table[5421] = 14'b0000101_0110100;
		logarithm_table[5422] = 14'b0000101_0110100;
		logarithm_table[5423] = 14'b0000101_0110100;
		logarithm_table[5424] = 14'b0000101_0110100;
		logarithm_table[5425] = 14'b0000101_0110100;
		logarithm_table[5426] = 14'b0000101_0110100;
		logarithm_table[5427] = 14'b0000101_0110100;
		logarithm_table[5428] = 14'b0000101_0110100;
		logarithm_table[5429] = 14'b0000101_0110100;
		logarithm_table[5430] = 14'b0000101_0110100;
		logarithm_table[5431] = 14'b0000101_0110100;
		logarithm_table[5432] = 14'b0000101_0110100;
		logarithm_table[5433] = 14'b0000101_0110100;
		logarithm_table[5434] = 14'b0000101_0110100;
		logarithm_table[5435] = 14'b0000101_0110100;
		logarithm_table[5436] = 14'b0000101_0110100;
		logarithm_table[5437] = 14'b0000101_0110100;
		logarithm_table[5438] = 14'b0000101_0110100;
		logarithm_table[5439] = 14'b0000101_0110100;
		logarithm_table[5440] = 14'b0000101_0110100;
		logarithm_table[5441] = 14'b0000101_0110100;
		logarithm_table[5442] = 14'b0000101_0110100;
		logarithm_table[5443] = 14'b0000101_0110101;
		logarithm_table[5444] = 14'b0000101_0110101;
		logarithm_table[5445] = 14'b0000101_0110101;
		logarithm_table[5446] = 14'b0000101_0110101;
		logarithm_table[5447] = 14'b0000101_0110101;
		logarithm_table[5448] = 14'b0000101_0110101;
		logarithm_table[5449] = 14'b0000101_0110101;
		logarithm_table[5450] = 14'b0000101_0110101;
		logarithm_table[5451] = 14'b0000101_0110101;
		logarithm_table[5452] = 14'b0000101_0110101;
		logarithm_table[5453] = 14'b0000101_0110101;
		logarithm_table[5454] = 14'b0000101_0110101;
		logarithm_table[5455] = 14'b0000101_0110101;
		logarithm_table[5456] = 14'b0000101_0110101;
		logarithm_table[5457] = 14'b0000101_0110101;
		logarithm_table[5458] = 14'b0000101_0110101;
		logarithm_table[5459] = 14'b0000101_0110101;
		logarithm_table[5460] = 14'b0000101_0110101;
		logarithm_table[5461] = 14'b0000101_0110101;
		logarithm_table[5462] = 14'b0000101_0110101;
		logarithm_table[5463] = 14'b0000101_0110101;
		logarithm_table[5464] = 14'b0000101_0110101;
		logarithm_table[5465] = 14'b0000101_0110101;
		logarithm_table[5466] = 14'b0000101_0110101;
		logarithm_table[5467] = 14'b0000101_0110101;
		logarithm_table[5468] = 14'b0000101_0110101;
		logarithm_table[5469] = 14'b0000101_0110101;
		logarithm_table[5470] = 14'b0000101_0110101;
		logarithm_table[5471] = 14'b0000101_0110101;
		logarithm_table[5472] = 14'b0000101_0110101;
		logarithm_table[5473] = 14'b0000101_0110110;
		logarithm_table[5474] = 14'b0000101_0110110;
		logarithm_table[5475] = 14'b0000101_0110110;
		logarithm_table[5476] = 14'b0000101_0110110;
		logarithm_table[5477] = 14'b0000101_0110110;
		logarithm_table[5478] = 14'b0000101_0110110;
		logarithm_table[5479] = 14'b0000101_0110110;
		logarithm_table[5480] = 14'b0000101_0110110;
		logarithm_table[5481] = 14'b0000101_0110110;
		logarithm_table[5482] = 14'b0000101_0110110;
		logarithm_table[5483] = 14'b0000101_0110110;
		logarithm_table[5484] = 14'b0000101_0110110;
		logarithm_table[5485] = 14'b0000101_0110110;
		logarithm_table[5486] = 14'b0000101_0110110;
		logarithm_table[5487] = 14'b0000101_0110110;
		logarithm_table[5488] = 14'b0000101_0110110;
		logarithm_table[5489] = 14'b0000101_0110110;
		logarithm_table[5490] = 14'b0000101_0110110;
		logarithm_table[5491] = 14'b0000101_0110110;
		logarithm_table[5492] = 14'b0000101_0110110;
		logarithm_table[5493] = 14'b0000101_0110110;
		logarithm_table[5494] = 14'b0000101_0110110;
		logarithm_table[5495] = 14'b0000101_0110110;
		logarithm_table[5496] = 14'b0000101_0110110;
		logarithm_table[5497] = 14'b0000101_0110110;
		logarithm_table[5498] = 14'b0000101_0110110;
		logarithm_table[5499] = 14'b0000101_0110110;
		logarithm_table[5500] = 14'b0000101_0110110;
		logarithm_table[5501] = 14'b0000101_0110110;
		logarithm_table[5502] = 14'b0000101_0110110;
		logarithm_table[5503] = 14'b0000101_0110111;
		logarithm_table[5504] = 14'b0000101_0110111;
		logarithm_table[5505] = 14'b0000101_0110111;
		logarithm_table[5506] = 14'b0000101_0110111;
		logarithm_table[5507] = 14'b0000101_0110111;
		logarithm_table[5508] = 14'b0000101_0110111;
		logarithm_table[5509] = 14'b0000101_0110111;
		logarithm_table[5510] = 14'b0000101_0110111;
		logarithm_table[5511] = 14'b0000101_0110111;
		logarithm_table[5512] = 14'b0000101_0110111;
		logarithm_table[5513] = 14'b0000101_0110111;
		logarithm_table[5514] = 14'b0000101_0110111;
		logarithm_table[5515] = 14'b0000101_0110111;
		logarithm_table[5516] = 14'b0000101_0110111;
		logarithm_table[5517] = 14'b0000101_0110111;
		logarithm_table[5518] = 14'b0000101_0110111;
		logarithm_table[5519] = 14'b0000101_0110111;
		logarithm_table[5520] = 14'b0000101_0110111;
		logarithm_table[5521] = 14'b0000101_0110111;
		logarithm_table[5522] = 14'b0000101_0110111;
		logarithm_table[5523] = 14'b0000101_0110111;
		logarithm_table[5524] = 14'b0000101_0110111;
		logarithm_table[5525] = 14'b0000101_0110111;
		logarithm_table[5526] = 14'b0000101_0110111;
		logarithm_table[5527] = 14'b0000101_0110111;
		logarithm_table[5528] = 14'b0000101_0110111;
		logarithm_table[5529] = 14'b0000101_0110111;
		logarithm_table[5530] = 14'b0000101_0110111;
		logarithm_table[5531] = 14'b0000101_0110111;
		logarithm_table[5532] = 14'b0000101_0110111;
		logarithm_table[5533] = 14'b0000101_0111000;
		logarithm_table[5534] = 14'b0000101_0111000;
		logarithm_table[5535] = 14'b0000101_0111000;
		logarithm_table[5536] = 14'b0000101_0111000;
		logarithm_table[5537] = 14'b0000101_0111000;
		logarithm_table[5538] = 14'b0000101_0111000;
		logarithm_table[5539] = 14'b0000101_0111000;
		logarithm_table[5540] = 14'b0000101_0111000;
		logarithm_table[5541] = 14'b0000101_0111000;
		logarithm_table[5542] = 14'b0000101_0111000;
		logarithm_table[5543] = 14'b0000101_0111000;
		logarithm_table[5544] = 14'b0000101_0111000;
		logarithm_table[5545] = 14'b0000101_0111000;
		logarithm_table[5546] = 14'b0000101_0111000;
		logarithm_table[5547] = 14'b0000101_0111000;
		logarithm_table[5548] = 14'b0000101_0111000;
		logarithm_table[5549] = 14'b0000101_0111000;
		logarithm_table[5550] = 14'b0000101_0111000;
		logarithm_table[5551] = 14'b0000101_0111000;
		logarithm_table[5552] = 14'b0000101_0111000;
		logarithm_table[5553] = 14'b0000101_0111000;
		logarithm_table[5554] = 14'b0000101_0111000;
		logarithm_table[5555] = 14'b0000101_0111000;
		logarithm_table[5556] = 14'b0000101_0111000;
		logarithm_table[5557] = 14'b0000101_0111000;
		logarithm_table[5558] = 14'b0000101_0111000;
		logarithm_table[5559] = 14'b0000101_0111000;
		logarithm_table[5560] = 14'b0000101_0111000;
		logarithm_table[5561] = 14'b0000101_0111000;
		logarithm_table[5562] = 14'b0000101_0111000;
		logarithm_table[5563] = 14'b0000101_0111001;
		logarithm_table[5564] = 14'b0000101_0111001;
		logarithm_table[5565] = 14'b0000101_0111001;
		logarithm_table[5566] = 14'b0000101_0111001;
		logarithm_table[5567] = 14'b0000101_0111001;
		logarithm_table[5568] = 14'b0000101_0111001;
		logarithm_table[5569] = 14'b0000101_0111001;
		logarithm_table[5570] = 14'b0000101_0111001;
		logarithm_table[5571] = 14'b0000101_0111001;
		logarithm_table[5572] = 14'b0000101_0111001;
		logarithm_table[5573] = 14'b0000101_0111001;
		logarithm_table[5574] = 14'b0000101_0111001;
		logarithm_table[5575] = 14'b0000101_0111001;
		logarithm_table[5576] = 14'b0000101_0111001;
		logarithm_table[5577] = 14'b0000101_0111001;
		logarithm_table[5578] = 14'b0000101_0111001;
		logarithm_table[5579] = 14'b0000101_0111001;
		logarithm_table[5580] = 14'b0000101_0111001;
		logarithm_table[5581] = 14'b0000101_0111001;
		logarithm_table[5582] = 14'b0000101_0111001;
		logarithm_table[5583] = 14'b0000101_0111001;
		logarithm_table[5584] = 14'b0000101_0111001;
		logarithm_table[5585] = 14'b0000101_0111001;
		logarithm_table[5586] = 14'b0000101_0111001;
		logarithm_table[5587] = 14'b0000101_0111001;
		logarithm_table[5588] = 14'b0000101_0111001;
		logarithm_table[5589] = 14'b0000101_0111001;
		logarithm_table[5590] = 14'b0000101_0111001;
		logarithm_table[5591] = 14'b0000101_0111001;
		logarithm_table[5592] = 14'b0000101_0111001;
		logarithm_table[5593] = 14'b0000101_0111010;
		logarithm_table[5594] = 14'b0000101_0111010;
		logarithm_table[5595] = 14'b0000101_0111010;
		logarithm_table[5596] = 14'b0000101_0111010;
		logarithm_table[5597] = 14'b0000101_0111010;
		logarithm_table[5598] = 14'b0000101_0111010;
		logarithm_table[5599] = 14'b0000101_0111010;
		logarithm_table[5600] = 14'b0000101_0111010;
		logarithm_table[5601] = 14'b0000101_0111010;
		logarithm_table[5602] = 14'b0000101_0111010;
		logarithm_table[5603] = 14'b0000101_0111010;
		logarithm_table[5604] = 14'b0000101_0111010;
		logarithm_table[5605] = 14'b0000101_0111010;
		logarithm_table[5606] = 14'b0000101_0111010;
		logarithm_table[5607] = 14'b0000101_0111010;
		logarithm_table[5608] = 14'b0000101_0111010;
		logarithm_table[5609] = 14'b0000101_0111010;
		logarithm_table[5610] = 14'b0000101_0111010;
		logarithm_table[5611] = 14'b0000101_0111010;
		logarithm_table[5612] = 14'b0000101_0111010;
		logarithm_table[5613] = 14'b0000101_0111010;
		logarithm_table[5614] = 14'b0000101_0111010;
		logarithm_table[5615] = 14'b0000101_0111010;
		logarithm_table[5616] = 14'b0000101_0111010;
		logarithm_table[5617] = 14'b0000101_0111010;
		logarithm_table[5618] = 14'b0000101_0111010;
		logarithm_table[5619] = 14'b0000101_0111010;
		logarithm_table[5620] = 14'b0000101_0111010;
		logarithm_table[5621] = 14'b0000101_0111010;
		logarithm_table[5622] = 14'b0000101_0111010;
		logarithm_table[5623] = 14'b0000101_0111011;
		logarithm_table[5624] = 14'b0000101_0111011;
		logarithm_table[5625] = 14'b0000101_0111011;
		logarithm_table[5626] = 14'b0000101_0111011;
		logarithm_table[5627] = 14'b0000101_0111011;
		logarithm_table[5628] = 14'b0000101_0111011;
		logarithm_table[5629] = 14'b0000101_0111011;
		logarithm_table[5630] = 14'b0000101_0111011;
		logarithm_table[5631] = 14'b0000101_0111011;
		logarithm_table[5632] = 14'b0000101_0111011;
		logarithm_table[5633] = 14'b0000101_0111011;
		logarithm_table[5634] = 14'b0000101_0111011;
		logarithm_table[5635] = 14'b0000101_0111011;
		logarithm_table[5636] = 14'b0000101_0111011;
		logarithm_table[5637] = 14'b0000101_0111011;
		logarithm_table[5638] = 14'b0000101_0111011;
		logarithm_table[5639] = 14'b0000101_0111011;
		logarithm_table[5640] = 14'b0000101_0111011;
		logarithm_table[5641] = 14'b0000101_0111011;
		logarithm_table[5642] = 14'b0000101_0111011;
		logarithm_table[5643] = 14'b0000101_0111011;
		logarithm_table[5644] = 14'b0000101_0111011;
		logarithm_table[5645] = 14'b0000101_0111011;
		logarithm_table[5646] = 14'b0000101_0111011;
		logarithm_table[5647] = 14'b0000101_0111011;
		logarithm_table[5648] = 14'b0000101_0111011;
		logarithm_table[5649] = 14'b0000101_0111011;
		logarithm_table[5650] = 14'b0000101_0111011;
		logarithm_table[5651] = 14'b0000101_0111011;
		logarithm_table[5652] = 14'b0000101_0111011;
		logarithm_table[5653] = 14'b0000101_0111011;
		logarithm_table[5654] = 14'b0000101_0111100;
		logarithm_table[5655] = 14'b0000101_0111100;
		logarithm_table[5656] = 14'b0000101_0111100;
		logarithm_table[5657] = 14'b0000101_0111100;
		logarithm_table[5658] = 14'b0000101_0111100;
		logarithm_table[5659] = 14'b0000101_0111100;
		logarithm_table[5660] = 14'b0000101_0111100;
		logarithm_table[5661] = 14'b0000101_0111100;
		logarithm_table[5662] = 14'b0000101_0111100;
		logarithm_table[5663] = 14'b0000101_0111100;
		logarithm_table[5664] = 14'b0000101_0111100;
		logarithm_table[5665] = 14'b0000101_0111100;
		logarithm_table[5666] = 14'b0000101_0111100;
		logarithm_table[5667] = 14'b0000101_0111100;
		logarithm_table[5668] = 14'b0000101_0111100;
		logarithm_table[5669] = 14'b0000101_0111100;
		logarithm_table[5670] = 14'b0000101_0111100;
		logarithm_table[5671] = 14'b0000101_0111100;
		logarithm_table[5672] = 14'b0000101_0111100;
		logarithm_table[5673] = 14'b0000101_0111100;
		logarithm_table[5674] = 14'b0000101_0111100;
		logarithm_table[5675] = 14'b0000101_0111100;
		logarithm_table[5676] = 14'b0000101_0111100;
		logarithm_table[5677] = 14'b0000101_0111100;
		logarithm_table[5678] = 14'b0000101_0111100;
		logarithm_table[5679] = 14'b0000101_0111100;
		logarithm_table[5680] = 14'b0000101_0111100;
		logarithm_table[5681] = 14'b0000101_0111100;
		logarithm_table[5682] = 14'b0000101_0111100;
		logarithm_table[5683] = 14'b0000101_0111100;
		logarithm_table[5684] = 14'b0000101_0111101;
		logarithm_table[5685] = 14'b0000101_0111101;
		logarithm_table[5686] = 14'b0000101_0111101;
		logarithm_table[5687] = 14'b0000101_0111101;
		logarithm_table[5688] = 14'b0000101_0111101;
		logarithm_table[5689] = 14'b0000101_0111101;
		logarithm_table[5690] = 14'b0000101_0111101;
		logarithm_table[5691] = 14'b0000101_0111101;
		logarithm_table[5692] = 14'b0000101_0111101;
		logarithm_table[5693] = 14'b0000101_0111101;
		logarithm_table[5694] = 14'b0000101_0111101;
		logarithm_table[5695] = 14'b0000101_0111101;
		logarithm_table[5696] = 14'b0000101_0111101;
		logarithm_table[5697] = 14'b0000101_0111101;
		logarithm_table[5698] = 14'b0000101_0111101;
		logarithm_table[5699] = 14'b0000101_0111101;
		logarithm_table[5700] = 14'b0000101_0111101;
		logarithm_table[5701] = 14'b0000101_0111101;
		logarithm_table[5702] = 14'b0000101_0111101;
		logarithm_table[5703] = 14'b0000101_0111101;
		logarithm_table[5704] = 14'b0000101_0111101;
		logarithm_table[5705] = 14'b0000101_0111101;
		logarithm_table[5706] = 14'b0000101_0111101;
		logarithm_table[5707] = 14'b0000101_0111101;
		logarithm_table[5708] = 14'b0000101_0111101;
		logarithm_table[5709] = 14'b0000101_0111101;
		logarithm_table[5710] = 14'b0000101_0111101;
		logarithm_table[5711] = 14'b0000101_0111101;
		logarithm_table[5712] = 14'b0000101_0111101;
		logarithm_table[5713] = 14'b0000101_0111101;
		logarithm_table[5714] = 14'b0000101_0111101;
		logarithm_table[5715] = 14'b0000101_0111110;
		logarithm_table[5716] = 14'b0000101_0111110;
		logarithm_table[5717] = 14'b0000101_0111110;
		logarithm_table[5718] = 14'b0000101_0111110;
		logarithm_table[5719] = 14'b0000101_0111110;
		logarithm_table[5720] = 14'b0000101_0111110;
		logarithm_table[5721] = 14'b0000101_0111110;
		logarithm_table[5722] = 14'b0000101_0111110;
		logarithm_table[5723] = 14'b0000101_0111110;
		logarithm_table[5724] = 14'b0000101_0111110;
		logarithm_table[5725] = 14'b0000101_0111110;
		logarithm_table[5726] = 14'b0000101_0111110;
		logarithm_table[5727] = 14'b0000101_0111110;
		logarithm_table[5728] = 14'b0000101_0111110;
		logarithm_table[5729] = 14'b0000101_0111110;
		logarithm_table[5730] = 14'b0000101_0111110;
		logarithm_table[5731] = 14'b0000101_0111110;
		logarithm_table[5732] = 14'b0000101_0111110;
		logarithm_table[5733] = 14'b0000101_0111110;
		logarithm_table[5734] = 14'b0000101_0111110;
		logarithm_table[5735] = 14'b0000101_0111110;
		logarithm_table[5736] = 14'b0000101_0111110;
		logarithm_table[5737] = 14'b0000101_0111110;
		logarithm_table[5738] = 14'b0000101_0111110;
		logarithm_table[5739] = 14'b0000101_0111110;
		logarithm_table[5740] = 14'b0000101_0111110;
		logarithm_table[5741] = 14'b0000101_0111110;
		logarithm_table[5742] = 14'b0000101_0111110;
		logarithm_table[5743] = 14'b0000101_0111110;
		logarithm_table[5744] = 14'b0000101_0111110;
		logarithm_table[5745] = 14'b0000101_0111110;
		logarithm_table[5746] = 14'b0000101_0111111;
		logarithm_table[5747] = 14'b0000101_0111111;
		logarithm_table[5748] = 14'b0000101_0111111;
		logarithm_table[5749] = 14'b0000101_0111111;
		logarithm_table[5750] = 14'b0000101_0111111;
		logarithm_table[5751] = 14'b0000101_0111111;
		logarithm_table[5752] = 14'b0000101_0111111;
		logarithm_table[5753] = 14'b0000101_0111111;
		logarithm_table[5754] = 14'b0000101_0111111;
		logarithm_table[5755] = 14'b0000101_0111111;
		logarithm_table[5756] = 14'b0000101_0111111;
		logarithm_table[5757] = 14'b0000101_0111111;
		logarithm_table[5758] = 14'b0000101_0111111;
		logarithm_table[5759] = 14'b0000101_0111111;
		logarithm_table[5760] = 14'b0000101_0111111;
		logarithm_table[5761] = 14'b0000101_0111111;
		logarithm_table[5762] = 14'b0000101_0111111;
		logarithm_table[5763] = 14'b0000101_0111111;
		logarithm_table[5764] = 14'b0000101_0111111;
		logarithm_table[5765] = 14'b0000101_0111111;
		logarithm_table[5766] = 14'b0000101_0111111;
		logarithm_table[5767] = 14'b0000101_0111111;
		logarithm_table[5768] = 14'b0000101_0111111;
		logarithm_table[5769] = 14'b0000101_0111111;
		logarithm_table[5770] = 14'b0000101_0111111;
		logarithm_table[5771] = 14'b0000101_0111111;
		logarithm_table[5772] = 14'b0000101_0111111;
		logarithm_table[5773] = 14'b0000101_0111111;
		logarithm_table[5774] = 14'b0000101_0111111;
		logarithm_table[5775] = 14'b0000101_0111111;
		logarithm_table[5776] = 14'b0000101_0111111;
		logarithm_table[5777] = 14'b0000101_1000000;
		logarithm_table[5778] = 14'b0000101_1000000;
		logarithm_table[5779] = 14'b0000101_1000000;
		logarithm_table[5780] = 14'b0000101_1000000;
		logarithm_table[5781] = 14'b0000101_1000000;
		logarithm_table[5782] = 14'b0000101_1000000;
		logarithm_table[5783] = 14'b0000101_1000000;
		logarithm_table[5784] = 14'b0000101_1000000;
		logarithm_table[5785] = 14'b0000101_1000000;
		logarithm_table[5786] = 14'b0000101_1000000;
		logarithm_table[5787] = 14'b0000101_1000000;
		logarithm_table[5788] = 14'b0000101_1000000;
		logarithm_table[5789] = 14'b0000101_1000000;
		logarithm_table[5790] = 14'b0000101_1000000;
		logarithm_table[5791] = 14'b0000101_1000000;
		logarithm_table[5792] = 14'b0000101_1000000;
		logarithm_table[5793] = 14'b0000101_1000000;
		logarithm_table[5794] = 14'b0000101_1000000;
		logarithm_table[5795] = 14'b0000101_1000000;
		logarithm_table[5796] = 14'b0000101_1000000;
		logarithm_table[5797] = 14'b0000101_1000000;
		logarithm_table[5798] = 14'b0000101_1000000;
		logarithm_table[5799] = 14'b0000101_1000000;
		logarithm_table[5800] = 14'b0000101_1000000;
		logarithm_table[5801] = 14'b0000101_1000000;
		logarithm_table[5802] = 14'b0000101_1000000;
		logarithm_table[5803] = 14'b0000101_1000000;
		logarithm_table[5804] = 14'b0000101_1000000;
		logarithm_table[5805] = 14'b0000101_1000000;
		logarithm_table[5806] = 14'b0000101_1000000;
		logarithm_table[5807] = 14'b0000101_1000000;
		logarithm_table[5808] = 14'b0000101_1000000;
		logarithm_table[5809] = 14'b0000101_1000001;
		logarithm_table[5810] = 14'b0000101_1000001;
		logarithm_table[5811] = 14'b0000101_1000001;
		logarithm_table[5812] = 14'b0000101_1000001;
		logarithm_table[5813] = 14'b0000101_1000001;
		logarithm_table[5814] = 14'b0000101_1000001;
		logarithm_table[5815] = 14'b0000101_1000001;
		logarithm_table[5816] = 14'b0000101_1000001;
		logarithm_table[5817] = 14'b0000101_1000001;
		logarithm_table[5818] = 14'b0000101_1000001;
		logarithm_table[5819] = 14'b0000101_1000001;
		logarithm_table[5820] = 14'b0000101_1000001;
		logarithm_table[5821] = 14'b0000101_1000001;
		logarithm_table[5822] = 14'b0000101_1000001;
		logarithm_table[5823] = 14'b0000101_1000001;
		logarithm_table[5824] = 14'b0000101_1000001;
		logarithm_table[5825] = 14'b0000101_1000001;
		logarithm_table[5826] = 14'b0000101_1000001;
		logarithm_table[5827] = 14'b0000101_1000001;
		logarithm_table[5828] = 14'b0000101_1000001;
		logarithm_table[5829] = 14'b0000101_1000001;
		logarithm_table[5830] = 14'b0000101_1000001;
		logarithm_table[5831] = 14'b0000101_1000001;
		logarithm_table[5832] = 14'b0000101_1000001;
		logarithm_table[5833] = 14'b0000101_1000001;
		logarithm_table[5834] = 14'b0000101_1000001;
		logarithm_table[5835] = 14'b0000101_1000001;
		logarithm_table[5836] = 14'b0000101_1000001;
		logarithm_table[5837] = 14'b0000101_1000001;
		logarithm_table[5838] = 14'b0000101_1000001;
		logarithm_table[5839] = 14'b0000101_1000001;
		logarithm_table[5840] = 14'b0000101_1000010;
		logarithm_table[5841] = 14'b0000101_1000010;
		logarithm_table[5842] = 14'b0000101_1000010;
		logarithm_table[5843] = 14'b0000101_1000010;
		logarithm_table[5844] = 14'b0000101_1000010;
		logarithm_table[5845] = 14'b0000101_1000010;
		logarithm_table[5846] = 14'b0000101_1000010;
		logarithm_table[5847] = 14'b0000101_1000010;
		logarithm_table[5848] = 14'b0000101_1000010;
		logarithm_table[5849] = 14'b0000101_1000010;
		logarithm_table[5850] = 14'b0000101_1000010;
		logarithm_table[5851] = 14'b0000101_1000010;
		logarithm_table[5852] = 14'b0000101_1000010;
		logarithm_table[5853] = 14'b0000101_1000010;
		logarithm_table[5854] = 14'b0000101_1000010;
		logarithm_table[5855] = 14'b0000101_1000010;
		logarithm_table[5856] = 14'b0000101_1000010;
		logarithm_table[5857] = 14'b0000101_1000010;
		logarithm_table[5858] = 14'b0000101_1000010;
		logarithm_table[5859] = 14'b0000101_1000010;
		logarithm_table[5860] = 14'b0000101_1000010;
		logarithm_table[5861] = 14'b0000101_1000010;
		logarithm_table[5862] = 14'b0000101_1000010;
		logarithm_table[5863] = 14'b0000101_1000010;
		logarithm_table[5864] = 14'b0000101_1000010;
		logarithm_table[5865] = 14'b0000101_1000010;
		logarithm_table[5866] = 14'b0000101_1000010;
		logarithm_table[5867] = 14'b0000101_1000010;
		logarithm_table[5868] = 14'b0000101_1000010;
		logarithm_table[5869] = 14'b0000101_1000010;
		logarithm_table[5870] = 14'b0000101_1000010;
		logarithm_table[5871] = 14'b0000101_1000010;
		logarithm_table[5872] = 14'b0000101_1000011;
		logarithm_table[5873] = 14'b0000101_1000011;
		logarithm_table[5874] = 14'b0000101_1000011;
		logarithm_table[5875] = 14'b0000101_1000011;
		logarithm_table[5876] = 14'b0000101_1000011;
		logarithm_table[5877] = 14'b0000101_1000011;
		logarithm_table[5878] = 14'b0000101_1000011;
		logarithm_table[5879] = 14'b0000101_1000011;
		logarithm_table[5880] = 14'b0000101_1000011;
		logarithm_table[5881] = 14'b0000101_1000011;
		logarithm_table[5882] = 14'b0000101_1000011;
		logarithm_table[5883] = 14'b0000101_1000011;
		logarithm_table[5884] = 14'b0000101_1000011;
		logarithm_table[5885] = 14'b0000101_1000011;
		logarithm_table[5886] = 14'b0000101_1000011;
		logarithm_table[5887] = 14'b0000101_1000011;
		logarithm_table[5888] = 14'b0000101_1000011;
		logarithm_table[5889] = 14'b0000101_1000011;
		logarithm_table[5890] = 14'b0000101_1000011;
		logarithm_table[5891] = 14'b0000101_1000011;
		logarithm_table[5892] = 14'b0000101_1000011;
		logarithm_table[5893] = 14'b0000101_1000011;
		logarithm_table[5894] = 14'b0000101_1000011;
		logarithm_table[5895] = 14'b0000101_1000011;
		logarithm_table[5896] = 14'b0000101_1000011;
		logarithm_table[5897] = 14'b0000101_1000011;
		logarithm_table[5898] = 14'b0000101_1000011;
		logarithm_table[5899] = 14'b0000101_1000011;
		logarithm_table[5900] = 14'b0000101_1000011;
		logarithm_table[5901] = 14'b0000101_1000011;
		logarithm_table[5902] = 14'b0000101_1000011;
		logarithm_table[5903] = 14'b0000101_1000011;
		logarithm_table[5904] = 14'b0000101_1000100;
		logarithm_table[5905] = 14'b0000101_1000100;
		logarithm_table[5906] = 14'b0000101_1000100;
		logarithm_table[5907] = 14'b0000101_1000100;
		logarithm_table[5908] = 14'b0000101_1000100;
		logarithm_table[5909] = 14'b0000101_1000100;
		logarithm_table[5910] = 14'b0000101_1000100;
		logarithm_table[5911] = 14'b0000101_1000100;
		logarithm_table[5912] = 14'b0000101_1000100;
		logarithm_table[5913] = 14'b0000101_1000100;
		logarithm_table[5914] = 14'b0000101_1000100;
		logarithm_table[5915] = 14'b0000101_1000100;
		logarithm_table[5916] = 14'b0000101_1000100;
		logarithm_table[5917] = 14'b0000101_1000100;
		logarithm_table[5918] = 14'b0000101_1000100;
		logarithm_table[5919] = 14'b0000101_1000100;
		logarithm_table[5920] = 14'b0000101_1000100;
		logarithm_table[5921] = 14'b0000101_1000100;
		logarithm_table[5922] = 14'b0000101_1000100;
		logarithm_table[5923] = 14'b0000101_1000100;
		logarithm_table[5924] = 14'b0000101_1000100;
		logarithm_table[5925] = 14'b0000101_1000100;
		logarithm_table[5926] = 14'b0000101_1000100;
		logarithm_table[5927] = 14'b0000101_1000100;
		logarithm_table[5928] = 14'b0000101_1000100;
		logarithm_table[5929] = 14'b0000101_1000100;
		logarithm_table[5930] = 14'b0000101_1000100;
		logarithm_table[5931] = 14'b0000101_1000100;
		logarithm_table[5932] = 14'b0000101_1000100;
		logarithm_table[5933] = 14'b0000101_1000100;
		logarithm_table[5934] = 14'b0000101_1000100;
		logarithm_table[5935] = 14'b0000101_1000100;
		logarithm_table[5936] = 14'b0000101_1000101;
		logarithm_table[5937] = 14'b0000101_1000101;
		logarithm_table[5938] = 14'b0000101_1000101;
		logarithm_table[5939] = 14'b0000101_1000101;
		logarithm_table[5940] = 14'b0000101_1000101;
		logarithm_table[5941] = 14'b0000101_1000101;
		logarithm_table[5942] = 14'b0000101_1000101;
		logarithm_table[5943] = 14'b0000101_1000101;
		logarithm_table[5944] = 14'b0000101_1000101;
		logarithm_table[5945] = 14'b0000101_1000101;
		logarithm_table[5946] = 14'b0000101_1000101;
		logarithm_table[5947] = 14'b0000101_1000101;
		logarithm_table[5948] = 14'b0000101_1000101;
		logarithm_table[5949] = 14'b0000101_1000101;
		logarithm_table[5950] = 14'b0000101_1000101;
		logarithm_table[5951] = 14'b0000101_1000101;
		logarithm_table[5952] = 14'b0000101_1000101;
		logarithm_table[5953] = 14'b0000101_1000101;
		logarithm_table[5954] = 14'b0000101_1000101;
		logarithm_table[5955] = 14'b0000101_1000101;
		logarithm_table[5956] = 14'b0000101_1000101;
		logarithm_table[5957] = 14'b0000101_1000101;
		logarithm_table[5958] = 14'b0000101_1000101;
		logarithm_table[5959] = 14'b0000101_1000101;
		logarithm_table[5960] = 14'b0000101_1000101;
		logarithm_table[5961] = 14'b0000101_1000101;
		logarithm_table[5962] = 14'b0000101_1000101;
		logarithm_table[5963] = 14'b0000101_1000101;
		logarithm_table[5964] = 14'b0000101_1000101;
		logarithm_table[5965] = 14'b0000101_1000101;
		logarithm_table[5966] = 14'b0000101_1000101;
		logarithm_table[5967] = 14'b0000101_1000101;
		logarithm_table[5968] = 14'b0000101_1000110;
		logarithm_table[5969] = 14'b0000101_1000110;
		logarithm_table[5970] = 14'b0000101_1000110;
		logarithm_table[5971] = 14'b0000101_1000110;
		logarithm_table[5972] = 14'b0000101_1000110;
		logarithm_table[5973] = 14'b0000101_1000110;
		logarithm_table[5974] = 14'b0000101_1000110;
		logarithm_table[5975] = 14'b0000101_1000110;
		logarithm_table[5976] = 14'b0000101_1000110;
		logarithm_table[5977] = 14'b0000101_1000110;
		logarithm_table[5978] = 14'b0000101_1000110;
		logarithm_table[5979] = 14'b0000101_1000110;
		logarithm_table[5980] = 14'b0000101_1000110;
		logarithm_table[5981] = 14'b0000101_1000110;
		logarithm_table[5982] = 14'b0000101_1000110;
		logarithm_table[5983] = 14'b0000101_1000110;
		logarithm_table[5984] = 14'b0000101_1000110;
		logarithm_table[5985] = 14'b0000101_1000110;
		logarithm_table[5986] = 14'b0000101_1000110;
		logarithm_table[5987] = 14'b0000101_1000110;
		logarithm_table[5988] = 14'b0000101_1000110;
		logarithm_table[5989] = 14'b0000101_1000110;
		logarithm_table[5990] = 14'b0000101_1000110;
		logarithm_table[5991] = 14'b0000101_1000110;
		logarithm_table[5992] = 14'b0000101_1000110;
		logarithm_table[5993] = 14'b0000101_1000110;
		logarithm_table[5994] = 14'b0000101_1000110;
		logarithm_table[5995] = 14'b0000101_1000110;
		logarithm_table[5996] = 14'b0000101_1000110;
		logarithm_table[5997] = 14'b0000101_1000110;
		logarithm_table[5998] = 14'b0000101_1000110;
		logarithm_table[5999] = 14'b0000101_1000110;
		logarithm_table[6000] = 14'b0000101_1000110;
		logarithm_table[6001] = 14'b0000101_1000111;
		logarithm_table[6002] = 14'b0000101_1000111;
		logarithm_table[6003] = 14'b0000101_1000111;
		logarithm_table[6004] = 14'b0000101_1000111;
		logarithm_table[6005] = 14'b0000101_1000111;
		logarithm_table[6006] = 14'b0000101_1000111;
		logarithm_table[6007] = 14'b0000101_1000111;
		logarithm_table[6008] = 14'b0000101_1000111;
		logarithm_table[6009] = 14'b0000101_1000111;
		logarithm_table[6010] = 14'b0000101_1000111;
		logarithm_table[6011] = 14'b0000101_1000111;
		logarithm_table[6012] = 14'b0000101_1000111;
		logarithm_table[6013] = 14'b0000101_1000111;
		logarithm_table[6014] = 14'b0000101_1000111;
		logarithm_table[6015] = 14'b0000101_1000111;
		logarithm_table[6016] = 14'b0000101_1000111;
		logarithm_table[6017] = 14'b0000101_1000111;
		logarithm_table[6018] = 14'b0000101_1000111;
		logarithm_table[6019] = 14'b0000101_1000111;
		logarithm_table[6020] = 14'b0000101_1000111;
		logarithm_table[6021] = 14'b0000101_1000111;
		logarithm_table[6022] = 14'b0000101_1000111;
		logarithm_table[6023] = 14'b0000101_1000111;
		logarithm_table[6024] = 14'b0000101_1000111;
		logarithm_table[6025] = 14'b0000101_1000111;
		logarithm_table[6026] = 14'b0000101_1000111;
		logarithm_table[6027] = 14'b0000101_1000111;
		logarithm_table[6028] = 14'b0000101_1000111;
		logarithm_table[6029] = 14'b0000101_1000111;
		logarithm_table[6030] = 14'b0000101_1000111;
		logarithm_table[6031] = 14'b0000101_1000111;
		logarithm_table[6032] = 14'b0000101_1000111;
		logarithm_table[6033] = 14'b0000101_1001000;
		logarithm_table[6034] = 14'b0000101_1001000;
		logarithm_table[6035] = 14'b0000101_1001000;
		logarithm_table[6036] = 14'b0000101_1001000;
		logarithm_table[6037] = 14'b0000101_1001000;
		logarithm_table[6038] = 14'b0000101_1001000;
		logarithm_table[6039] = 14'b0000101_1001000;
		logarithm_table[6040] = 14'b0000101_1001000;
		logarithm_table[6041] = 14'b0000101_1001000;
		logarithm_table[6042] = 14'b0000101_1001000;
		logarithm_table[6043] = 14'b0000101_1001000;
		logarithm_table[6044] = 14'b0000101_1001000;
		logarithm_table[6045] = 14'b0000101_1001000;
		logarithm_table[6046] = 14'b0000101_1001000;
		logarithm_table[6047] = 14'b0000101_1001000;
		logarithm_table[6048] = 14'b0000101_1001000;
		logarithm_table[6049] = 14'b0000101_1001000;
		logarithm_table[6050] = 14'b0000101_1001000;
		logarithm_table[6051] = 14'b0000101_1001000;
		logarithm_table[6052] = 14'b0000101_1001000;
		logarithm_table[6053] = 14'b0000101_1001000;
		logarithm_table[6054] = 14'b0000101_1001000;
		logarithm_table[6055] = 14'b0000101_1001000;
		logarithm_table[6056] = 14'b0000101_1001000;
		logarithm_table[6057] = 14'b0000101_1001000;
		logarithm_table[6058] = 14'b0000101_1001000;
		logarithm_table[6059] = 14'b0000101_1001000;
		logarithm_table[6060] = 14'b0000101_1001000;
		logarithm_table[6061] = 14'b0000101_1001000;
		logarithm_table[6062] = 14'b0000101_1001000;
		logarithm_table[6063] = 14'b0000101_1001000;
		logarithm_table[6064] = 14'b0000101_1001000;
		logarithm_table[6065] = 14'b0000101_1001000;
		logarithm_table[6066] = 14'b0000101_1001001;
		logarithm_table[6067] = 14'b0000101_1001001;
		logarithm_table[6068] = 14'b0000101_1001001;
		logarithm_table[6069] = 14'b0000101_1001001;
		logarithm_table[6070] = 14'b0000101_1001001;
		logarithm_table[6071] = 14'b0000101_1001001;
		logarithm_table[6072] = 14'b0000101_1001001;
		logarithm_table[6073] = 14'b0000101_1001001;
		logarithm_table[6074] = 14'b0000101_1001001;
		logarithm_table[6075] = 14'b0000101_1001001;
		logarithm_table[6076] = 14'b0000101_1001001;
		logarithm_table[6077] = 14'b0000101_1001001;
		logarithm_table[6078] = 14'b0000101_1001001;
		logarithm_table[6079] = 14'b0000101_1001001;
		logarithm_table[6080] = 14'b0000101_1001001;
		logarithm_table[6081] = 14'b0000101_1001001;
		logarithm_table[6082] = 14'b0000101_1001001;
		logarithm_table[6083] = 14'b0000101_1001001;
		logarithm_table[6084] = 14'b0000101_1001001;
		logarithm_table[6085] = 14'b0000101_1001001;
		logarithm_table[6086] = 14'b0000101_1001001;
		logarithm_table[6087] = 14'b0000101_1001001;
		logarithm_table[6088] = 14'b0000101_1001001;
		logarithm_table[6089] = 14'b0000101_1001001;
		logarithm_table[6090] = 14'b0000101_1001001;
		logarithm_table[6091] = 14'b0000101_1001001;
		logarithm_table[6092] = 14'b0000101_1001001;
		logarithm_table[6093] = 14'b0000101_1001001;
		logarithm_table[6094] = 14'b0000101_1001001;
		logarithm_table[6095] = 14'b0000101_1001001;
		logarithm_table[6096] = 14'b0000101_1001001;
		logarithm_table[6097] = 14'b0000101_1001001;
		logarithm_table[6098] = 14'b0000101_1001001;
		logarithm_table[6099] = 14'b0000101_1001010;
		logarithm_table[6100] = 14'b0000101_1001010;
		logarithm_table[6101] = 14'b0000101_1001010;
		logarithm_table[6102] = 14'b0000101_1001010;
		logarithm_table[6103] = 14'b0000101_1001010;
		logarithm_table[6104] = 14'b0000101_1001010;
		logarithm_table[6105] = 14'b0000101_1001010;
		logarithm_table[6106] = 14'b0000101_1001010;
		logarithm_table[6107] = 14'b0000101_1001010;
		logarithm_table[6108] = 14'b0000101_1001010;
		logarithm_table[6109] = 14'b0000101_1001010;
		logarithm_table[6110] = 14'b0000101_1001010;
		logarithm_table[6111] = 14'b0000101_1001010;
		logarithm_table[6112] = 14'b0000101_1001010;
		logarithm_table[6113] = 14'b0000101_1001010;
		logarithm_table[6114] = 14'b0000101_1001010;
		logarithm_table[6115] = 14'b0000101_1001010;
		logarithm_table[6116] = 14'b0000101_1001010;
		logarithm_table[6117] = 14'b0000101_1001010;
		logarithm_table[6118] = 14'b0000101_1001010;
		logarithm_table[6119] = 14'b0000101_1001010;
		logarithm_table[6120] = 14'b0000101_1001010;
		logarithm_table[6121] = 14'b0000101_1001010;
		logarithm_table[6122] = 14'b0000101_1001010;
		logarithm_table[6123] = 14'b0000101_1001010;
		logarithm_table[6124] = 14'b0000101_1001010;
		logarithm_table[6125] = 14'b0000101_1001010;
		logarithm_table[6126] = 14'b0000101_1001010;
		logarithm_table[6127] = 14'b0000101_1001010;
		logarithm_table[6128] = 14'b0000101_1001010;
		logarithm_table[6129] = 14'b0000101_1001010;
		logarithm_table[6130] = 14'b0000101_1001010;
		logarithm_table[6131] = 14'b0000101_1001010;
		logarithm_table[6132] = 14'b0000101_1001011;
		logarithm_table[6133] = 14'b0000101_1001011;
		logarithm_table[6134] = 14'b0000101_1001011;
		logarithm_table[6135] = 14'b0000101_1001011;
		logarithm_table[6136] = 14'b0000101_1001011;
		logarithm_table[6137] = 14'b0000101_1001011;
		logarithm_table[6138] = 14'b0000101_1001011;
		logarithm_table[6139] = 14'b0000101_1001011;
		logarithm_table[6140] = 14'b0000101_1001011;
		logarithm_table[6141] = 14'b0000101_1001011;
		logarithm_table[6142] = 14'b0000101_1001011;
		logarithm_table[6143] = 14'b0000101_1001011;
		logarithm_table[6144] = 14'b0000101_1001011;
		logarithm_table[6145] = 14'b0000101_1001011;
		logarithm_table[6146] = 14'b0000101_1001011;
		logarithm_table[6147] = 14'b0000101_1001011;
		logarithm_table[6148] = 14'b0000101_1001011;
		logarithm_table[6149] = 14'b0000101_1001011;
		logarithm_table[6150] = 14'b0000101_1001011;
		logarithm_table[6151] = 14'b0000101_1001011;
		logarithm_table[6152] = 14'b0000101_1001011;
		logarithm_table[6153] = 14'b0000101_1001011;
		logarithm_table[6154] = 14'b0000101_1001011;
		logarithm_table[6155] = 14'b0000101_1001011;
		logarithm_table[6156] = 14'b0000101_1001011;
		logarithm_table[6157] = 14'b0000101_1001011;
		logarithm_table[6158] = 14'b0000101_1001011;
		logarithm_table[6159] = 14'b0000101_1001011;
		logarithm_table[6160] = 14'b0000101_1001011;
		logarithm_table[6161] = 14'b0000101_1001011;
		logarithm_table[6162] = 14'b0000101_1001011;
		logarithm_table[6163] = 14'b0000101_1001011;
		logarithm_table[6164] = 14'b0000101_1001011;
		logarithm_table[6165] = 14'b0000101_1001100;
		logarithm_table[6166] = 14'b0000101_1001100;
		logarithm_table[6167] = 14'b0000101_1001100;
		logarithm_table[6168] = 14'b0000101_1001100;
		logarithm_table[6169] = 14'b0000101_1001100;
		logarithm_table[6170] = 14'b0000101_1001100;
		logarithm_table[6171] = 14'b0000101_1001100;
		logarithm_table[6172] = 14'b0000101_1001100;
		logarithm_table[6173] = 14'b0000101_1001100;
		logarithm_table[6174] = 14'b0000101_1001100;
		logarithm_table[6175] = 14'b0000101_1001100;
		logarithm_table[6176] = 14'b0000101_1001100;
		logarithm_table[6177] = 14'b0000101_1001100;
		logarithm_table[6178] = 14'b0000101_1001100;
		logarithm_table[6179] = 14'b0000101_1001100;
		logarithm_table[6180] = 14'b0000101_1001100;
		logarithm_table[6181] = 14'b0000101_1001100;
		logarithm_table[6182] = 14'b0000101_1001100;
		logarithm_table[6183] = 14'b0000101_1001100;
		logarithm_table[6184] = 14'b0000101_1001100;
		logarithm_table[6185] = 14'b0000101_1001100;
		logarithm_table[6186] = 14'b0000101_1001100;
		logarithm_table[6187] = 14'b0000101_1001100;
		logarithm_table[6188] = 14'b0000101_1001100;
		logarithm_table[6189] = 14'b0000101_1001100;
		logarithm_table[6190] = 14'b0000101_1001100;
		logarithm_table[6191] = 14'b0000101_1001100;
		logarithm_table[6192] = 14'b0000101_1001100;
		logarithm_table[6193] = 14'b0000101_1001100;
		logarithm_table[6194] = 14'b0000101_1001100;
		logarithm_table[6195] = 14'b0000101_1001100;
		logarithm_table[6196] = 14'b0000101_1001100;
		logarithm_table[6197] = 14'b0000101_1001100;
		logarithm_table[6198] = 14'b0000101_1001100;
		logarithm_table[6199] = 14'b0000101_1001101;
		logarithm_table[6200] = 14'b0000101_1001101;
		logarithm_table[6201] = 14'b0000101_1001101;
		logarithm_table[6202] = 14'b0000101_1001101;
		logarithm_table[6203] = 14'b0000101_1001101;
		logarithm_table[6204] = 14'b0000101_1001101;
		logarithm_table[6205] = 14'b0000101_1001101;
		logarithm_table[6206] = 14'b0000101_1001101;
		logarithm_table[6207] = 14'b0000101_1001101;
		logarithm_table[6208] = 14'b0000101_1001101;
		logarithm_table[6209] = 14'b0000101_1001101;
		logarithm_table[6210] = 14'b0000101_1001101;
		logarithm_table[6211] = 14'b0000101_1001101;
		logarithm_table[6212] = 14'b0000101_1001101;
		logarithm_table[6213] = 14'b0000101_1001101;
		logarithm_table[6214] = 14'b0000101_1001101;
		logarithm_table[6215] = 14'b0000101_1001101;
		logarithm_table[6216] = 14'b0000101_1001101;
		logarithm_table[6217] = 14'b0000101_1001101;
		logarithm_table[6218] = 14'b0000101_1001101;
		logarithm_table[6219] = 14'b0000101_1001101;
		logarithm_table[6220] = 14'b0000101_1001101;
		logarithm_table[6221] = 14'b0000101_1001101;
		logarithm_table[6222] = 14'b0000101_1001101;
		logarithm_table[6223] = 14'b0000101_1001101;
		logarithm_table[6224] = 14'b0000101_1001101;
		logarithm_table[6225] = 14'b0000101_1001101;
		logarithm_table[6226] = 14'b0000101_1001101;
		logarithm_table[6227] = 14'b0000101_1001101;
		logarithm_table[6228] = 14'b0000101_1001101;
		logarithm_table[6229] = 14'b0000101_1001101;
		logarithm_table[6230] = 14'b0000101_1001101;
		logarithm_table[6231] = 14'b0000101_1001101;
		logarithm_table[6232] = 14'b0000101_1001110;
		logarithm_table[6233] = 14'b0000101_1001110;
		logarithm_table[6234] = 14'b0000101_1001110;
		logarithm_table[6235] = 14'b0000101_1001110;
		logarithm_table[6236] = 14'b0000101_1001110;
		logarithm_table[6237] = 14'b0000101_1001110;
		logarithm_table[6238] = 14'b0000101_1001110;
		logarithm_table[6239] = 14'b0000101_1001110;
		logarithm_table[6240] = 14'b0000101_1001110;
		logarithm_table[6241] = 14'b0000101_1001110;
		logarithm_table[6242] = 14'b0000101_1001110;
		logarithm_table[6243] = 14'b0000101_1001110;
		logarithm_table[6244] = 14'b0000101_1001110;
		logarithm_table[6245] = 14'b0000101_1001110;
		logarithm_table[6246] = 14'b0000101_1001110;
		logarithm_table[6247] = 14'b0000101_1001110;
		logarithm_table[6248] = 14'b0000101_1001110;
		logarithm_table[6249] = 14'b0000101_1001110;
		logarithm_table[6250] = 14'b0000101_1001110;
		logarithm_table[6251] = 14'b0000101_1001110;
		logarithm_table[6252] = 14'b0000101_1001110;
		logarithm_table[6253] = 14'b0000101_1001110;
		logarithm_table[6254] = 14'b0000101_1001110;
		logarithm_table[6255] = 14'b0000101_1001110;
		logarithm_table[6256] = 14'b0000101_1001110;
		logarithm_table[6257] = 14'b0000101_1001110;
		logarithm_table[6258] = 14'b0000101_1001110;
		logarithm_table[6259] = 14'b0000101_1001110;
		logarithm_table[6260] = 14'b0000101_1001110;
		logarithm_table[6261] = 14'b0000101_1001110;
		logarithm_table[6262] = 14'b0000101_1001110;
		logarithm_table[6263] = 14'b0000101_1001110;
		logarithm_table[6264] = 14'b0000101_1001110;
		logarithm_table[6265] = 14'b0000101_1001110;
		logarithm_table[6266] = 14'b0000101_1001111;
		logarithm_table[6267] = 14'b0000101_1001111;
		logarithm_table[6268] = 14'b0000101_1001111;
		logarithm_table[6269] = 14'b0000101_1001111;
		logarithm_table[6270] = 14'b0000101_1001111;
		logarithm_table[6271] = 14'b0000101_1001111;
		logarithm_table[6272] = 14'b0000101_1001111;
		logarithm_table[6273] = 14'b0000101_1001111;
		logarithm_table[6274] = 14'b0000101_1001111;
		logarithm_table[6275] = 14'b0000101_1001111;
		logarithm_table[6276] = 14'b0000101_1001111;
		logarithm_table[6277] = 14'b0000101_1001111;
		logarithm_table[6278] = 14'b0000101_1001111;
		logarithm_table[6279] = 14'b0000101_1001111;
		logarithm_table[6280] = 14'b0000101_1001111;
		logarithm_table[6281] = 14'b0000101_1001111;
		logarithm_table[6282] = 14'b0000101_1001111;
		logarithm_table[6283] = 14'b0000101_1001111;
		logarithm_table[6284] = 14'b0000101_1001111;
		logarithm_table[6285] = 14'b0000101_1001111;
		logarithm_table[6286] = 14'b0000101_1001111;
		logarithm_table[6287] = 14'b0000101_1001111;
		logarithm_table[6288] = 14'b0000101_1001111;
		logarithm_table[6289] = 14'b0000101_1001111;
		logarithm_table[6290] = 14'b0000101_1001111;
		logarithm_table[6291] = 14'b0000101_1001111;
		logarithm_table[6292] = 14'b0000101_1001111;
		logarithm_table[6293] = 14'b0000101_1001111;
		logarithm_table[6294] = 14'b0000101_1001111;
		logarithm_table[6295] = 14'b0000101_1001111;
		logarithm_table[6296] = 14'b0000101_1001111;
		logarithm_table[6297] = 14'b0000101_1001111;
		logarithm_table[6298] = 14'b0000101_1001111;
		logarithm_table[6299] = 14'b0000101_1001111;
		logarithm_table[6300] = 14'b0000101_1010000;
		logarithm_table[6301] = 14'b0000101_1010000;
		logarithm_table[6302] = 14'b0000101_1010000;
		logarithm_table[6303] = 14'b0000101_1010000;
		logarithm_table[6304] = 14'b0000101_1010000;
		logarithm_table[6305] = 14'b0000101_1010000;
		logarithm_table[6306] = 14'b0000101_1010000;
		logarithm_table[6307] = 14'b0000101_1010000;
		logarithm_table[6308] = 14'b0000101_1010000;
		logarithm_table[6309] = 14'b0000101_1010000;
		logarithm_table[6310] = 14'b0000101_1010000;
		logarithm_table[6311] = 14'b0000101_1010000;
		logarithm_table[6312] = 14'b0000101_1010000;
		logarithm_table[6313] = 14'b0000101_1010000;
		logarithm_table[6314] = 14'b0000101_1010000;
		logarithm_table[6315] = 14'b0000101_1010000;
		logarithm_table[6316] = 14'b0000101_1010000;
		logarithm_table[6317] = 14'b0000101_1010000;
		logarithm_table[6318] = 14'b0000101_1010000;
		logarithm_table[6319] = 14'b0000101_1010000;
		logarithm_table[6320] = 14'b0000101_1010000;
		logarithm_table[6321] = 14'b0000101_1010000;
		logarithm_table[6322] = 14'b0000101_1010000;
		logarithm_table[6323] = 14'b0000101_1010000;
		logarithm_table[6324] = 14'b0000101_1010000;
		logarithm_table[6325] = 14'b0000101_1010000;
		logarithm_table[6326] = 14'b0000101_1010000;
		logarithm_table[6327] = 14'b0000101_1010000;
		logarithm_table[6328] = 14'b0000101_1010000;
		logarithm_table[6329] = 14'b0000101_1010000;
		logarithm_table[6330] = 14'b0000101_1010000;
		logarithm_table[6331] = 14'b0000101_1010000;
		logarithm_table[6332] = 14'b0000101_1010000;
		logarithm_table[6333] = 14'b0000101_1010000;
		logarithm_table[6334] = 14'b0000101_1010000;
		logarithm_table[6335] = 14'b0000101_1010001;
		logarithm_table[6336] = 14'b0000101_1010001;
		logarithm_table[6337] = 14'b0000101_1010001;
		logarithm_table[6338] = 14'b0000101_1010001;
		logarithm_table[6339] = 14'b0000101_1010001;
		logarithm_table[6340] = 14'b0000101_1010001;
		logarithm_table[6341] = 14'b0000101_1010001;
		logarithm_table[6342] = 14'b0000101_1010001;
		logarithm_table[6343] = 14'b0000101_1010001;
		logarithm_table[6344] = 14'b0000101_1010001;
		logarithm_table[6345] = 14'b0000101_1010001;
		logarithm_table[6346] = 14'b0000101_1010001;
		logarithm_table[6347] = 14'b0000101_1010001;
		logarithm_table[6348] = 14'b0000101_1010001;
		logarithm_table[6349] = 14'b0000101_1010001;
		logarithm_table[6350] = 14'b0000101_1010001;
		logarithm_table[6351] = 14'b0000101_1010001;
		logarithm_table[6352] = 14'b0000101_1010001;
		logarithm_table[6353] = 14'b0000101_1010001;
		logarithm_table[6354] = 14'b0000101_1010001;
		logarithm_table[6355] = 14'b0000101_1010001;
		logarithm_table[6356] = 14'b0000101_1010001;
		logarithm_table[6357] = 14'b0000101_1010001;
		logarithm_table[6358] = 14'b0000101_1010001;
		logarithm_table[6359] = 14'b0000101_1010001;
		logarithm_table[6360] = 14'b0000101_1010001;
		logarithm_table[6361] = 14'b0000101_1010001;
		logarithm_table[6362] = 14'b0000101_1010001;
		logarithm_table[6363] = 14'b0000101_1010001;
		logarithm_table[6364] = 14'b0000101_1010001;
		logarithm_table[6365] = 14'b0000101_1010001;
		logarithm_table[6366] = 14'b0000101_1010001;
		logarithm_table[6367] = 14'b0000101_1010001;
		logarithm_table[6368] = 14'b0000101_1010001;
		logarithm_table[6369] = 14'b0000101_1010010;
		logarithm_table[6370] = 14'b0000101_1010010;
		logarithm_table[6371] = 14'b0000101_1010010;
		logarithm_table[6372] = 14'b0000101_1010010;
		logarithm_table[6373] = 14'b0000101_1010010;
		logarithm_table[6374] = 14'b0000101_1010010;
		logarithm_table[6375] = 14'b0000101_1010010;
		logarithm_table[6376] = 14'b0000101_1010010;
		logarithm_table[6377] = 14'b0000101_1010010;
		logarithm_table[6378] = 14'b0000101_1010010;
		logarithm_table[6379] = 14'b0000101_1010010;
		logarithm_table[6380] = 14'b0000101_1010010;
		logarithm_table[6381] = 14'b0000101_1010010;
		logarithm_table[6382] = 14'b0000101_1010010;
		logarithm_table[6383] = 14'b0000101_1010010;
		logarithm_table[6384] = 14'b0000101_1010010;
		logarithm_table[6385] = 14'b0000101_1010010;
		logarithm_table[6386] = 14'b0000101_1010010;
		logarithm_table[6387] = 14'b0000101_1010010;
		logarithm_table[6388] = 14'b0000101_1010010;
		logarithm_table[6389] = 14'b0000101_1010010;
		logarithm_table[6390] = 14'b0000101_1010010;
		logarithm_table[6391] = 14'b0000101_1010010;
		logarithm_table[6392] = 14'b0000101_1010010;
		logarithm_table[6393] = 14'b0000101_1010010;
		logarithm_table[6394] = 14'b0000101_1010010;
		logarithm_table[6395] = 14'b0000101_1010010;
		logarithm_table[6396] = 14'b0000101_1010010;
		logarithm_table[6397] = 14'b0000101_1010010;
		logarithm_table[6398] = 14'b0000101_1010010;
		logarithm_table[6399] = 14'b0000101_1010010;
		logarithm_table[6400] = 14'b0000101_1010010;
		logarithm_table[6401] = 14'b0000101_1010010;
		logarithm_table[6402] = 14'b0000101_1010010;
		logarithm_table[6403] = 14'b0000101_1010011;
		logarithm_table[6404] = 14'b0000101_1010011;
		logarithm_table[6405] = 14'b0000101_1010011;
		logarithm_table[6406] = 14'b0000101_1010011;
		logarithm_table[6407] = 14'b0000101_1010011;
		logarithm_table[6408] = 14'b0000101_1010011;
		logarithm_table[6409] = 14'b0000101_1010011;
		logarithm_table[6410] = 14'b0000101_1010011;
		logarithm_table[6411] = 14'b0000101_1010011;
		logarithm_table[6412] = 14'b0000101_1010011;
		logarithm_table[6413] = 14'b0000101_1010011;
		logarithm_table[6414] = 14'b0000101_1010011;
		logarithm_table[6415] = 14'b0000101_1010011;
		logarithm_table[6416] = 14'b0000101_1010011;
		logarithm_table[6417] = 14'b0000101_1010011;
		logarithm_table[6418] = 14'b0000101_1010011;
		logarithm_table[6419] = 14'b0000101_1010011;
		logarithm_table[6420] = 14'b0000101_1010011;
		logarithm_table[6421] = 14'b0000101_1010011;
		logarithm_table[6422] = 14'b0000101_1010011;
		logarithm_table[6423] = 14'b0000101_1010011;
		logarithm_table[6424] = 14'b0000101_1010011;
		logarithm_table[6425] = 14'b0000101_1010011;
		logarithm_table[6426] = 14'b0000101_1010011;
		logarithm_table[6427] = 14'b0000101_1010011;
		logarithm_table[6428] = 14'b0000101_1010011;
		logarithm_table[6429] = 14'b0000101_1010011;
		logarithm_table[6430] = 14'b0000101_1010011;
		logarithm_table[6431] = 14'b0000101_1010011;
		logarithm_table[6432] = 14'b0000101_1010011;
		logarithm_table[6433] = 14'b0000101_1010011;
		logarithm_table[6434] = 14'b0000101_1010011;
		logarithm_table[6435] = 14'b0000101_1010011;
		logarithm_table[6436] = 14'b0000101_1010011;
		logarithm_table[6437] = 14'b0000101_1010011;
		logarithm_table[6438] = 14'b0000101_1010100;
		logarithm_table[6439] = 14'b0000101_1010100;
		logarithm_table[6440] = 14'b0000101_1010100;
		logarithm_table[6441] = 14'b0000101_1010100;
		logarithm_table[6442] = 14'b0000101_1010100;
		logarithm_table[6443] = 14'b0000101_1010100;
		logarithm_table[6444] = 14'b0000101_1010100;
		logarithm_table[6445] = 14'b0000101_1010100;
		logarithm_table[6446] = 14'b0000101_1010100;
		logarithm_table[6447] = 14'b0000101_1010100;
		logarithm_table[6448] = 14'b0000101_1010100;
		logarithm_table[6449] = 14'b0000101_1010100;
		logarithm_table[6450] = 14'b0000101_1010100;
		logarithm_table[6451] = 14'b0000101_1010100;
		logarithm_table[6452] = 14'b0000101_1010100;
		logarithm_table[6453] = 14'b0000101_1010100;
		logarithm_table[6454] = 14'b0000101_1010100;
		logarithm_table[6455] = 14'b0000101_1010100;
		logarithm_table[6456] = 14'b0000101_1010100;
		logarithm_table[6457] = 14'b0000101_1010100;
		logarithm_table[6458] = 14'b0000101_1010100;
		logarithm_table[6459] = 14'b0000101_1010100;
		logarithm_table[6460] = 14'b0000101_1010100;
		logarithm_table[6461] = 14'b0000101_1010100;
		logarithm_table[6462] = 14'b0000101_1010100;
		logarithm_table[6463] = 14'b0000101_1010100;
		logarithm_table[6464] = 14'b0000101_1010100;
		logarithm_table[6465] = 14'b0000101_1010100;
		logarithm_table[6466] = 14'b0000101_1010100;
		logarithm_table[6467] = 14'b0000101_1010100;
		logarithm_table[6468] = 14'b0000101_1010100;
		logarithm_table[6469] = 14'b0000101_1010100;
		logarithm_table[6470] = 14'b0000101_1010100;
		logarithm_table[6471] = 14'b0000101_1010100;
		logarithm_table[6472] = 14'b0000101_1010100;
		logarithm_table[6473] = 14'b0000101_1010101;
		logarithm_table[6474] = 14'b0000101_1010101;
		logarithm_table[6475] = 14'b0000101_1010101;
		logarithm_table[6476] = 14'b0000101_1010101;
		logarithm_table[6477] = 14'b0000101_1010101;
		logarithm_table[6478] = 14'b0000101_1010101;
		logarithm_table[6479] = 14'b0000101_1010101;
		logarithm_table[6480] = 14'b0000101_1010101;
		logarithm_table[6481] = 14'b0000101_1010101;
		logarithm_table[6482] = 14'b0000101_1010101;
		logarithm_table[6483] = 14'b0000101_1010101;
		logarithm_table[6484] = 14'b0000101_1010101;
		logarithm_table[6485] = 14'b0000101_1010101;
		logarithm_table[6486] = 14'b0000101_1010101;
		logarithm_table[6487] = 14'b0000101_1010101;
		logarithm_table[6488] = 14'b0000101_1010101;
		logarithm_table[6489] = 14'b0000101_1010101;
		logarithm_table[6490] = 14'b0000101_1010101;
		logarithm_table[6491] = 14'b0000101_1010101;
		logarithm_table[6492] = 14'b0000101_1010101;
		logarithm_table[6493] = 14'b0000101_1010101;
		logarithm_table[6494] = 14'b0000101_1010101;
		logarithm_table[6495] = 14'b0000101_1010101;
		logarithm_table[6496] = 14'b0000101_1010101;
		logarithm_table[6497] = 14'b0000101_1010101;
		logarithm_table[6498] = 14'b0000101_1010101;
		logarithm_table[6499] = 14'b0000101_1010101;
		logarithm_table[6500] = 14'b0000101_1010101;
		logarithm_table[6501] = 14'b0000101_1010101;
		logarithm_table[6502] = 14'b0000101_1010101;
		logarithm_table[6503] = 14'b0000101_1010101;
		logarithm_table[6504] = 14'b0000101_1010101;
		logarithm_table[6505] = 14'b0000101_1010101;
		logarithm_table[6506] = 14'b0000101_1010101;
		logarithm_table[6507] = 14'b0000101_1010101;
		logarithm_table[6508] = 14'b0000101_1010110;
		logarithm_table[6509] = 14'b0000101_1010110;
		logarithm_table[6510] = 14'b0000101_1010110;
		logarithm_table[6511] = 14'b0000101_1010110;
		logarithm_table[6512] = 14'b0000101_1010110;
		logarithm_table[6513] = 14'b0000101_1010110;
		logarithm_table[6514] = 14'b0000101_1010110;
		logarithm_table[6515] = 14'b0000101_1010110;
		logarithm_table[6516] = 14'b0000101_1010110;
		logarithm_table[6517] = 14'b0000101_1010110;
		logarithm_table[6518] = 14'b0000101_1010110;
		logarithm_table[6519] = 14'b0000101_1010110;
		logarithm_table[6520] = 14'b0000101_1010110;
		logarithm_table[6521] = 14'b0000101_1010110;
		logarithm_table[6522] = 14'b0000101_1010110;
		logarithm_table[6523] = 14'b0000101_1010110;
		logarithm_table[6524] = 14'b0000101_1010110;
		logarithm_table[6525] = 14'b0000101_1010110;
		logarithm_table[6526] = 14'b0000101_1010110;
		logarithm_table[6527] = 14'b0000101_1010110;
		logarithm_table[6528] = 14'b0000101_1010110;
		logarithm_table[6529] = 14'b0000101_1010110;
		logarithm_table[6530] = 14'b0000101_1010110;
		logarithm_table[6531] = 14'b0000101_1010110;
		logarithm_table[6532] = 14'b0000101_1010110;
		logarithm_table[6533] = 14'b0000101_1010110;
		logarithm_table[6534] = 14'b0000101_1010110;
		logarithm_table[6535] = 14'b0000101_1010110;
		logarithm_table[6536] = 14'b0000101_1010110;
		logarithm_table[6537] = 14'b0000101_1010110;
		logarithm_table[6538] = 14'b0000101_1010110;
		logarithm_table[6539] = 14'b0000101_1010110;
		logarithm_table[6540] = 14'b0000101_1010110;
		logarithm_table[6541] = 14'b0000101_1010110;
		logarithm_table[6542] = 14'b0000101_1010110;
		logarithm_table[6543] = 14'b0000101_1010110;
		logarithm_table[6544] = 14'b0000101_1010111;
		logarithm_table[6545] = 14'b0000101_1010111;
		logarithm_table[6546] = 14'b0000101_1010111;
		logarithm_table[6547] = 14'b0000101_1010111;
		logarithm_table[6548] = 14'b0000101_1010111;
		logarithm_table[6549] = 14'b0000101_1010111;
		logarithm_table[6550] = 14'b0000101_1010111;
		logarithm_table[6551] = 14'b0000101_1010111;
		logarithm_table[6552] = 14'b0000101_1010111;
		logarithm_table[6553] = 14'b0000101_1010111;
		logarithm_table[6554] = 14'b0000101_1010111;
		logarithm_table[6555] = 14'b0000101_1010111;
		logarithm_table[6556] = 14'b0000101_1010111;
		logarithm_table[6557] = 14'b0000101_1010111;
		logarithm_table[6558] = 14'b0000101_1010111;
		logarithm_table[6559] = 14'b0000101_1010111;
		logarithm_table[6560] = 14'b0000101_1010111;
		logarithm_table[6561] = 14'b0000101_1010111;
		logarithm_table[6562] = 14'b0000101_1010111;
		logarithm_table[6563] = 14'b0000101_1010111;
		logarithm_table[6564] = 14'b0000101_1010111;
		logarithm_table[6565] = 14'b0000101_1010111;
		logarithm_table[6566] = 14'b0000101_1010111;
		logarithm_table[6567] = 14'b0000101_1010111;
		logarithm_table[6568] = 14'b0000101_1010111;
		logarithm_table[6569] = 14'b0000101_1010111;
		logarithm_table[6570] = 14'b0000101_1010111;
		logarithm_table[6571] = 14'b0000101_1010111;
		logarithm_table[6572] = 14'b0000101_1010111;
		logarithm_table[6573] = 14'b0000101_1010111;
		logarithm_table[6574] = 14'b0000101_1010111;
		logarithm_table[6575] = 14'b0000101_1010111;
		logarithm_table[6576] = 14'b0000101_1010111;
		logarithm_table[6577] = 14'b0000101_1010111;
		logarithm_table[6578] = 14'b0000101_1010111;
		logarithm_table[6579] = 14'b0000101_1011000;
		logarithm_table[6580] = 14'b0000101_1011000;
		logarithm_table[6581] = 14'b0000101_1011000;
		logarithm_table[6582] = 14'b0000101_1011000;
		logarithm_table[6583] = 14'b0000101_1011000;
		logarithm_table[6584] = 14'b0000101_1011000;
		logarithm_table[6585] = 14'b0000101_1011000;
		logarithm_table[6586] = 14'b0000101_1011000;
		logarithm_table[6587] = 14'b0000101_1011000;
		logarithm_table[6588] = 14'b0000101_1011000;
		logarithm_table[6589] = 14'b0000101_1011000;
		logarithm_table[6590] = 14'b0000101_1011000;
		logarithm_table[6591] = 14'b0000101_1011000;
		logarithm_table[6592] = 14'b0000101_1011000;
		logarithm_table[6593] = 14'b0000101_1011000;
		logarithm_table[6594] = 14'b0000101_1011000;
		logarithm_table[6595] = 14'b0000101_1011000;
		logarithm_table[6596] = 14'b0000101_1011000;
		logarithm_table[6597] = 14'b0000101_1011000;
		logarithm_table[6598] = 14'b0000101_1011000;
		logarithm_table[6599] = 14'b0000101_1011000;
		logarithm_table[6600] = 14'b0000101_1011000;
		logarithm_table[6601] = 14'b0000101_1011000;
		logarithm_table[6602] = 14'b0000101_1011000;
		logarithm_table[6603] = 14'b0000101_1011000;
		logarithm_table[6604] = 14'b0000101_1011000;
		logarithm_table[6605] = 14'b0000101_1011000;
		logarithm_table[6606] = 14'b0000101_1011000;
		logarithm_table[6607] = 14'b0000101_1011000;
		logarithm_table[6608] = 14'b0000101_1011000;
		logarithm_table[6609] = 14'b0000101_1011000;
		logarithm_table[6610] = 14'b0000101_1011000;
		logarithm_table[6611] = 14'b0000101_1011000;
		logarithm_table[6612] = 14'b0000101_1011000;
		logarithm_table[6613] = 14'b0000101_1011000;
		logarithm_table[6614] = 14'b0000101_1011000;
		logarithm_table[6615] = 14'b0000101_1011001;
		logarithm_table[6616] = 14'b0000101_1011001;
		logarithm_table[6617] = 14'b0000101_1011001;
		logarithm_table[6618] = 14'b0000101_1011001;
		logarithm_table[6619] = 14'b0000101_1011001;
		logarithm_table[6620] = 14'b0000101_1011001;
		logarithm_table[6621] = 14'b0000101_1011001;
		logarithm_table[6622] = 14'b0000101_1011001;
		logarithm_table[6623] = 14'b0000101_1011001;
		logarithm_table[6624] = 14'b0000101_1011001;
		logarithm_table[6625] = 14'b0000101_1011001;
		logarithm_table[6626] = 14'b0000101_1011001;
		logarithm_table[6627] = 14'b0000101_1011001;
		logarithm_table[6628] = 14'b0000101_1011001;
		logarithm_table[6629] = 14'b0000101_1011001;
		logarithm_table[6630] = 14'b0000101_1011001;
		logarithm_table[6631] = 14'b0000101_1011001;
		logarithm_table[6632] = 14'b0000101_1011001;
		logarithm_table[6633] = 14'b0000101_1011001;
		logarithm_table[6634] = 14'b0000101_1011001;
		logarithm_table[6635] = 14'b0000101_1011001;
		logarithm_table[6636] = 14'b0000101_1011001;
		logarithm_table[6637] = 14'b0000101_1011001;
		logarithm_table[6638] = 14'b0000101_1011001;
		logarithm_table[6639] = 14'b0000101_1011001;
		logarithm_table[6640] = 14'b0000101_1011001;
		logarithm_table[6641] = 14'b0000101_1011001;
		logarithm_table[6642] = 14'b0000101_1011001;
		logarithm_table[6643] = 14'b0000101_1011001;
		logarithm_table[6644] = 14'b0000101_1011001;
		logarithm_table[6645] = 14'b0000101_1011001;
		logarithm_table[6646] = 14'b0000101_1011001;
		logarithm_table[6647] = 14'b0000101_1011001;
		logarithm_table[6648] = 14'b0000101_1011001;
		logarithm_table[6649] = 14'b0000101_1011001;
		logarithm_table[6650] = 14'b0000101_1011001;
		logarithm_table[6651] = 14'b0000101_1011010;
		logarithm_table[6652] = 14'b0000101_1011010;
		logarithm_table[6653] = 14'b0000101_1011010;
		logarithm_table[6654] = 14'b0000101_1011010;
		logarithm_table[6655] = 14'b0000101_1011010;
		logarithm_table[6656] = 14'b0000101_1011010;
		logarithm_table[6657] = 14'b0000101_1011010;
		logarithm_table[6658] = 14'b0000101_1011010;
		logarithm_table[6659] = 14'b0000101_1011010;
		logarithm_table[6660] = 14'b0000101_1011010;
		logarithm_table[6661] = 14'b0000101_1011010;
		logarithm_table[6662] = 14'b0000101_1011010;
		logarithm_table[6663] = 14'b0000101_1011010;
		logarithm_table[6664] = 14'b0000101_1011010;
		logarithm_table[6665] = 14'b0000101_1011010;
		logarithm_table[6666] = 14'b0000101_1011010;
		logarithm_table[6667] = 14'b0000101_1011010;
		logarithm_table[6668] = 14'b0000101_1011010;
		logarithm_table[6669] = 14'b0000101_1011010;
		logarithm_table[6670] = 14'b0000101_1011010;
		logarithm_table[6671] = 14'b0000101_1011010;
		logarithm_table[6672] = 14'b0000101_1011010;
		logarithm_table[6673] = 14'b0000101_1011010;
		logarithm_table[6674] = 14'b0000101_1011010;
		logarithm_table[6675] = 14'b0000101_1011010;
		logarithm_table[6676] = 14'b0000101_1011010;
		logarithm_table[6677] = 14'b0000101_1011010;
		logarithm_table[6678] = 14'b0000101_1011010;
		logarithm_table[6679] = 14'b0000101_1011010;
		logarithm_table[6680] = 14'b0000101_1011010;
		logarithm_table[6681] = 14'b0000101_1011010;
		logarithm_table[6682] = 14'b0000101_1011010;
		logarithm_table[6683] = 14'b0000101_1011010;
		logarithm_table[6684] = 14'b0000101_1011010;
		logarithm_table[6685] = 14'b0000101_1011010;
		logarithm_table[6686] = 14'b0000101_1011010;
		logarithm_table[6687] = 14'b0000101_1011011;
		logarithm_table[6688] = 14'b0000101_1011011;
		logarithm_table[6689] = 14'b0000101_1011011;
		logarithm_table[6690] = 14'b0000101_1011011;
		logarithm_table[6691] = 14'b0000101_1011011;
		logarithm_table[6692] = 14'b0000101_1011011;
		logarithm_table[6693] = 14'b0000101_1011011;
		logarithm_table[6694] = 14'b0000101_1011011;
		logarithm_table[6695] = 14'b0000101_1011011;
		logarithm_table[6696] = 14'b0000101_1011011;
		logarithm_table[6697] = 14'b0000101_1011011;
		logarithm_table[6698] = 14'b0000101_1011011;
		logarithm_table[6699] = 14'b0000101_1011011;
		logarithm_table[6700] = 14'b0000101_1011011;
		logarithm_table[6701] = 14'b0000101_1011011;
		logarithm_table[6702] = 14'b0000101_1011011;
		logarithm_table[6703] = 14'b0000101_1011011;
		logarithm_table[6704] = 14'b0000101_1011011;
		logarithm_table[6705] = 14'b0000101_1011011;
		logarithm_table[6706] = 14'b0000101_1011011;
		logarithm_table[6707] = 14'b0000101_1011011;
		logarithm_table[6708] = 14'b0000101_1011011;
		logarithm_table[6709] = 14'b0000101_1011011;
		logarithm_table[6710] = 14'b0000101_1011011;
		logarithm_table[6711] = 14'b0000101_1011011;
		logarithm_table[6712] = 14'b0000101_1011011;
		logarithm_table[6713] = 14'b0000101_1011011;
		logarithm_table[6714] = 14'b0000101_1011011;
		logarithm_table[6715] = 14'b0000101_1011011;
		logarithm_table[6716] = 14'b0000101_1011011;
		logarithm_table[6717] = 14'b0000101_1011011;
		logarithm_table[6718] = 14'b0000101_1011011;
		logarithm_table[6719] = 14'b0000101_1011011;
		logarithm_table[6720] = 14'b0000101_1011011;
		logarithm_table[6721] = 14'b0000101_1011011;
		logarithm_table[6722] = 14'b0000101_1011011;
		logarithm_table[6723] = 14'b0000101_1011100;
		logarithm_table[6724] = 14'b0000101_1011100;
		logarithm_table[6725] = 14'b0000101_1011100;
		logarithm_table[6726] = 14'b0000101_1011100;
		logarithm_table[6727] = 14'b0000101_1011100;
		logarithm_table[6728] = 14'b0000101_1011100;
		logarithm_table[6729] = 14'b0000101_1011100;
		logarithm_table[6730] = 14'b0000101_1011100;
		logarithm_table[6731] = 14'b0000101_1011100;
		logarithm_table[6732] = 14'b0000101_1011100;
		logarithm_table[6733] = 14'b0000101_1011100;
		logarithm_table[6734] = 14'b0000101_1011100;
		logarithm_table[6735] = 14'b0000101_1011100;
		logarithm_table[6736] = 14'b0000101_1011100;
		logarithm_table[6737] = 14'b0000101_1011100;
		logarithm_table[6738] = 14'b0000101_1011100;
		logarithm_table[6739] = 14'b0000101_1011100;
		logarithm_table[6740] = 14'b0000101_1011100;
		logarithm_table[6741] = 14'b0000101_1011100;
		logarithm_table[6742] = 14'b0000101_1011100;
		logarithm_table[6743] = 14'b0000101_1011100;
		logarithm_table[6744] = 14'b0000101_1011100;
		logarithm_table[6745] = 14'b0000101_1011100;
		logarithm_table[6746] = 14'b0000101_1011100;
		logarithm_table[6747] = 14'b0000101_1011100;
		logarithm_table[6748] = 14'b0000101_1011100;
		logarithm_table[6749] = 14'b0000101_1011100;
		logarithm_table[6750] = 14'b0000101_1011100;
		logarithm_table[6751] = 14'b0000101_1011100;
		logarithm_table[6752] = 14'b0000101_1011100;
		logarithm_table[6753] = 14'b0000101_1011100;
		logarithm_table[6754] = 14'b0000101_1011100;
		logarithm_table[6755] = 14'b0000101_1011100;
		logarithm_table[6756] = 14'b0000101_1011100;
		logarithm_table[6757] = 14'b0000101_1011100;
		logarithm_table[6758] = 14'b0000101_1011100;
		logarithm_table[6759] = 14'b0000101_1011100;
		logarithm_table[6760] = 14'b0000101_1011101;
		logarithm_table[6761] = 14'b0000101_1011101;
		logarithm_table[6762] = 14'b0000101_1011101;
		logarithm_table[6763] = 14'b0000101_1011101;
		logarithm_table[6764] = 14'b0000101_1011101;
		logarithm_table[6765] = 14'b0000101_1011101;
		logarithm_table[6766] = 14'b0000101_1011101;
		logarithm_table[6767] = 14'b0000101_1011101;
		logarithm_table[6768] = 14'b0000101_1011101;
		logarithm_table[6769] = 14'b0000101_1011101;
		logarithm_table[6770] = 14'b0000101_1011101;
		logarithm_table[6771] = 14'b0000101_1011101;
		logarithm_table[6772] = 14'b0000101_1011101;
		logarithm_table[6773] = 14'b0000101_1011101;
		logarithm_table[6774] = 14'b0000101_1011101;
		logarithm_table[6775] = 14'b0000101_1011101;
		logarithm_table[6776] = 14'b0000101_1011101;
		logarithm_table[6777] = 14'b0000101_1011101;
		logarithm_table[6778] = 14'b0000101_1011101;
		logarithm_table[6779] = 14'b0000101_1011101;
		logarithm_table[6780] = 14'b0000101_1011101;
		logarithm_table[6781] = 14'b0000101_1011101;
		logarithm_table[6782] = 14'b0000101_1011101;
		logarithm_table[6783] = 14'b0000101_1011101;
		logarithm_table[6784] = 14'b0000101_1011101;
		logarithm_table[6785] = 14'b0000101_1011101;
		logarithm_table[6786] = 14'b0000101_1011101;
		logarithm_table[6787] = 14'b0000101_1011101;
		logarithm_table[6788] = 14'b0000101_1011101;
		logarithm_table[6789] = 14'b0000101_1011101;
		logarithm_table[6790] = 14'b0000101_1011101;
		logarithm_table[6791] = 14'b0000101_1011101;
		logarithm_table[6792] = 14'b0000101_1011101;
		logarithm_table[6793] = 14'b0000101_1011101;
		logarithm_table[6794] = 14'b0000101_1011101;
		logarithm_table[6795] = 14'b0000101_1011101;
		logarithm_table[6796] = 14'b0000101_1011110;
		logarithm_table[6797] = 14'b0000101_1011110;
		logarithm_table[6798] = 14'b0000101_1011110;
		logarithm_table[6799] = 14'b0000101_1011110;
		logarithm_table[6800] = 14'b0000101_1011110;
		logarithm_table[6801] = 14'b0000101_1011110;
		logarithm_table[6802] = 14'b0000101_1011110;
		logarithm_table[6803] = 14'b0000101_1011110;
		logarithm_table[6804] = 14'b0000101_1011110;
		logarithm_table[6805] = 14'b0000101_1011110;
		logarithm_table[6806] = 14'b0000101_1011110;
		logarithm_table[6807] = 14'b0000101_1011110;
		logarithm_table[6808] = 14'b0000101_1011110;
		logarithm_table[6809] = 14'b0000101_1011110;
		logarithm_table[6810] = 14'b0000101_1011110;
		logarithm_table[6811] = 14'b0000101_1011110;
		logarithm_table[6812] = 14'b0000101_1011110;
		logarithm_table[6813] = 14'b0000101_1011110;
		logarithm_table[6814] = 14'b0000101_1011110;
		logarithm_table[6815] = 14'b0000101_1011110;
		logarithm_table[6816] = 14'b0000101_1011110;
		logarithm_table[6817] = 14'b0000101_1011110;
		logarithm_table[6818] = 14'b0000101_1011110;
		logarithm_table[6819] = 14'b0000101_1011110;
		logarithm_table[6820] = 14'b0000101_1011110;
		logarithm_table[6821] = 14'b0000101_1011110;
		logarithm_table[6822] = 14'b0000101_1011110;
		logarithm_table[6823] = 14'b0000101_1011110;
		logarithm_table[6824] = 14'b0000101_1011110;
		logarithm_table[6825] = 14'b0000101_1011110;
		logarithm_table[6826] = 14'b0000101_1011110;
		logarithm_table[6827] = 14'b0000101_1011110;
		logarithm_table[6828] = 14'b0000101_1011110;
		logarithm_table[6829] = 14'b0000101_1011110;
		logarithm_table[6830] = 14'b0000101_1011110;
		logarithm_table[6831] = 14'b0000101_1011110;
		logarithm_table[6832] = 14'b0000101_1011110;
		logarithm_table[6833] = 14'b0000101_1011111;
		logarithm_table[6834] = 14'b0000101_1011111;
		logarithm_table[6835] = 14'b0000101_1011111;
		logarithm_table[6836] = 14'b0000101_1011111;
		logarithm_table[6837] = 14'b0000101_1011111;
		logarithm_table[6838] = 14'b0000101_1011111;
		logarithm_table[6839] = 14'b0000101_1011111;
		logarithm_table[6840] = 14'b0000101_1011111;
		logarithm_table[6841] = 14'b0000101_1011111;
		logarithm_table[6842] = 14'b0000101_1011111;
		logarithm_table[6843] = 14'b0000101_1011111;
		logarithm_table[6844] = 14'b0000101_1011111;
		logarithm_table[6845] = 14'b0000101_1011111;
		logarithm_table[6846] = 14'b0000101_1011111;
		logarithm_table[6847] = 14'b0000101_1011111;
		logarithm_table[6848] = 14'b0000101_1011111;
		logarithm_table[6849] = 14'b0000101_1011111;
		logarithm_table[6850] = 14'b0000101_1011111;
		logarithm_table[6851] = 14'b0000101_1011111;
		logarithm_table[6852] = 14'b0000101_1011111;
		logarithm_table[6853] = 14'b0000101_1011111;
		logarithm_table[6854] = 14'b0000101_1011111;
		logarithm_table[6855] = 14'b0000101_1011111;
		logarithm_table[6856] = 14'b0000101_1011111;
		logarithm_table[6857] = 14'b0000101_1011111;
		logarithm_table[6858] = 14'b0000101_1011111;
		logarithm_table[6859] = 14'b0000101_1011111;
		logarithm_table[6860] = 14'b0000101_1011111;
		logarithm_table[6861] = 14'b0000101_1011111;
		logarithm_table[6862] = 14'b0000101_1011111;
		logarithm_table[6863] = 14'b0000101_1011111;
		logarithm_table[6864] = 14'b0000101_1011111;
		logarithm_table[6865] = 14'b0000101_1011111;
		logarithm_table[6866] = 14'b0000101_1011111;
		logarithm_table[6867] = 14'b0000101_1011111;
		logarithm_table[6868] = 14'b0000101_1011111;
		logarithm_table[6869] = 14'b0000101_1011111;
		logarithm_table[6870] = 14'b0000101_1100000;
		logarithm_table[6871] = 14'b0000101_1100000;
		logarithm_table[6872] = 14'b0000101_1100000;
		logarithm_table[6873] = 14'b0000101_1100000;
		logarithm_table[6874] = 14'b0000101_1100000;
		logarithm_table[6875] = 14'b0000101_1100000;
		logarithm_table[6876] = 14'b0000101_1100000;
		logarithm_table[6877] = 14'b0000101_1100000;
		logarithm_table[6878] = 14'b0000101_1100000;
		logarithm_table[6879] = 14'b0000101_1100000;
		logarithm_table[6880] = 14'b0000101_1100000;
		logarithm_table[6881] = 14'b0000101_1100000;
		logarithm_table[6882] = 14'b0000101_1100000;
		logarithm_table[6883] = 14'b0000101_1100000;
		logarithm_table[6884] = 14'b0000101_1100000;
		logarithm_table[6885] = 14'b0000101_1100000;
		logarithm_table[6886] = 14'b0000101_1100000;
		logarithm_table[6887] = 14'b0000101_1100000;
		logarithm_table[6888] = 14'b0000101_1100000;
		logarithm_table[6889] = 14'b0000101_1100000;
		logarithm_table[6890] = 14'b0000101_1100000;
		logarithm_table[6891] = 14'b0000101_1100000;
		logarithm_table[6892] = 14'b0000101_1100000;
		logarithm_table[6893] = 14'b0000101_1100000;
		logarithm_table[6894] = 14'b0000101_1100000;
		logarithm_table[6895] = 14'b0000101_1100000;
		logarithm_table[6896] = 14'b0000101_1100000;
		logarithm_table[6897] = 14'b0000101_1100000;
		logarithm_table[6898] = 14'b0000101_1100000;
		logarithm_table[6899] = 14'b0000101_1100000;
		logarithm_table[6900] = 14'b0000101_1100000;
		logarithm_table[6901] = 14'b0000101_1100000;
		logarithm_table[6902] = 14'b0000101_1100000;
		logarithm_table[6903] = 14'b0000101_1100000;
		logarithm_table[6904] = 14'b0000101_1100000;
		logarithm_table[6905] = 14'b0000101_1100000;
		logarithm_table[6906] = 14'b0000101_1100000;
		logarithm_table[6907] = 14'b0000101_1100000;
		logarithm_table[6908] = 14'b0000101_1100001;
		logarithm_table[6909] = 14'b0000101_1100001;
		logarithm_table[6910] = 14'b0000101_1100001;
		logarithm_table[6911] = 14'b0000101_1100001;
		logarithm_table[6912] = 14'b0000101_1100001;
		logarithm_table[6913] = 14'b0000101_1100001;
		logarithm_table[6914] = 14'b0000101_1100001;
		logarithm_table[6915] = 14'b0000101_1100001;
		logarithm_table[6916] = 14'b0000101_1100001;
		logarithm_table[6917] = 14'b0000101_1100001;
		logarithm_table[6918] = 14'b0000101_1100001;
		logarithm_table[6919] = 14'b0000101_1100001;
		logarithm_table[6920] = 14'b0000101_1100001;
		logarithm_table[6921] = 14'b0000101_1100001;
		logarithm_table[6922] = 14'b0000101_1100001;
		logarithm_table[6923] = 14'b0000101_1100001;
		logarithm_table[6924] = 14'b0000101_1100001;
		logarithm_table[6925] = 14'b0000101_1100001;
		logarithm_table[6926] = 14'b0000101_1100001;
		logarithm_table[6927] = 14'b0000101_1100001;
		logarithm_table[6928] = 14'b0000101_1100001;
		logarithm_table[6929] = 14'b0000101_1100001;
		logarithm_table[6930] = 14'b0000101_1100001;
		logarithm_table[6931] = 14'b0000101_1100001;
		logarithm_table[6932] = 14'b0000101_1100001;
		logarithm_table[6933] = 14'b0000101_1100001;
		logarithm_table[6934] = 14'b0000101_1100001;
		logarithm_table[6935] = 14'b0000101_1100001;
		logarithm_table[6936] = 14'b0000101_1100001;
		logarithm_table[6937] = 14'b0000101_1100001;
		logarithm_table[6938] = 14'b0000101_1100001;
		logarithm_table[6939] = 14'b0000101_1100001;
		logarithm_table[6940] = 14'b0000101_1100001;
		logarithm_table[6941] = 14'b0000101_1100001;
		logarithm_table[6942] = 14'b0000101_1100001;
		logarithm_table[6943] = 14'b0000101_1100001;
		logarithm_table[6944] = 14'b0000101_1100001;
		logarithm_table[6945] = 14'b0000101_1100010;
		logarithm_table[6946] = 14'b0000101_1100010;
		logarithm_table[6947] = 14'b0000101_1100010;
		logarithm_table[6948] = 14'b0000101_1100010;
		logarithm_table[6949] = 14'b0000101_1100010;
		logarithm_table[6950] = 14'b0000101_1100010;
		logarithm_table[6951] = 14'b0000101_1100010;
		logarithm_table[6952] = 14'b0000101_1100010;
		logarithm_table[6953] = 14'b0000101_1100010;
		logarithm_table[6954] = 14'b0000101_1100010;
		logarithm_table[6955] = 14'b0000101_1100010;
		logarithm_table[6956] = 14'b0000101_1100010;
		logarithm_table[6957] = 14'b0000101_1100010;
		logarithm_table[6958] = 14'b0000101_1100010;
		logarithm_table[6959] = 14'b0000101_1100010;
		logarithm_table[6960] = 14'b0000101_1100010;
		logarithm_table[6961] = 14'b0000101_1100010;
		logarithm_table[6962] = 14'b0000101_1100010;
		logarithm_table[6963] = 14'b0000101_1100010;
		logarithm_table[6964] = 14'b0000101_1100010;
		logarithm_table[6965] = 14'b0000101_1100010;
		logarithm_table[6966] = 14'b0000101_1100010;
		logarithm_table[6967] = 14'b0000101_1100010;
		logarithm_table[6968] = 14'b0000101_1100010;
		logarithm_table[6969] = 14'b0000101_1100010;
		logarithm_table[6970] = 14'b0000101_1100010;
		logarithm_table[6971] = 14'b0000101_1100010;
		logarithm_table[6972] = 14'b0000101_1100010;
		logarithm_table[6973] = 14'b0000101_1100010;
		logarithm_table[6974] = 14'b0000101_1100010;
		logarithm_table[6975] = 14'b0000101_1100010;
		logarithm_table[6976] = 14'b0000101_1100010;
		logarithm_table[6977] = 14'b0000101_1100010;
		logarithm_table[6978] = 14'b0000101_1100010;
		logarithm_table[6979] = 14'b0000101_1100010;
		logarithm_table[6980] = 14'b0000101_1100010;
		logarithm_table[6981] = 14'b0000101_1100010;
		logarithm_table[6982] = 14'b0000101_1100010;
		logarithm_table[6983] = 14'b0000101_1100011;
		logarithm_table[6984] = 14'b0000101_1100011;
		logarithm_table[6985] = 14'b0000101_1100011;
		logarithm_table[6986] = 14'b0000101_1100011;
		logarithm_table[6987] = 14'b0000101_1100011;
		logarithm_table[6988] = 14'b0000101_1100011;
		logarithm_table[6989] = 14'b0000101_1100011;
		logarithm_table[6990] = 14'b0000101_1100011;
		logarithm_table[6991] = 14'b0000101_1100011;
		logarithm_table[6992] = 14'b0000101_1100011;
		logarithm_table[6993] = 14'b0000101_1100011;
		logarithm_table[6994] = 14'b0000101_1100011;
		logarithm_table[6995] = 14'b0000101_1100011;
		logarithm_table[6996] = 14'b0000101_1100011;
		logarithm_table[6997] = 14'b0000101_1100011;
		logarithm_table[6998] = 14'b0000101_1100011;
		logarithm_table[6999] = 14'b0000101_1100011;
		logarithm_table[7000] = 14'b0000101_1100011;
		logarithm_table[7001] = 14'b0000101_1100011;
		logarithm_table[7002] = 14'b0000101_1100011;
		logarithm_table[7003] = 14'b0000101_1100011;
		logarithm_table[7004] = 14'b0000101_1100011;
		logarithm_table[7005] = 14'b0000101_1100011;
		logarithm_table[7006] = 14'b0000101_1100011;
		logarithm_table[7007] = 14'b0000101_1100011;
		logarithm_table[7008] = 14'b0000101_1100011;
		logarithm_table[7009] = 14'b0000101_1100011;
		logarithm_table[7010] = 14'b0000101_1100011;
		logarithm_table[7011] = 14'b0000101_1100011;
		logarithm_table[7012] = 14'b0000101_1100011;
		logarithm_table[7013] = 14'b0000101_1100011;
		logarithm_table[7014] = 14'b0000101_1100011;
		logarithm_table[7015] = 14'b0000101_1100011;
		logarithm_table[7016] = 14'b0000101_1100011;
		logarithm_table[7017] = 14'b0000101_1100011;
		logarithm_table[7018] = 14'b0000101_1100011;
		logarithm_table[7019] = 14'b0000101_1100011;
		logarithm_table[7020] = 14'b0000101_1100011;
		logarithm_table[7021] = 14'b0000101_1100100;
		logarithm_table[7022] = 14'b0000101_1100100;
		logarithm_table[7023] = 14'b0000101_1100100;
		logarithm_table[7024] = 14'b0000101_1100100;
		logarithm_table[7025] = 14'b0000101_1100100;
		logarithm_table[7026] = 14'b0000101_1100100;
		logarithm_table[7027] = 14'b0000101_1100100;
		logarithm_table[7028] = 14'b0000101_1100100;
		logarithm_table[7029] = 14'b0000101_1100100;
		logarithm_table[7030] = 14'b0000101_1100100;
		logarithm_table[7031] = 14'b0000101_1100100;
		logarithm_table[7032] = 14'b0000101_1100100;
		logarithm_table[7033] = 14'b0000101_1100100;
		logarithm_table[7034] = 14'b0000101_1100100;
		logarithm_table[7035] = 14'b0000101_1100100;
		logarithm_table[7036] = 14'b0000101_1100100;
		logarithm_table[7037] = 14'b0000101_1100100;
		logarithm_table[7038] = 14'b0000101_1100100;
		logarithm_table[7039] = 14'b0000101_1100100;
		logarithm_table[7040] = 14'b0000101_1100100;
		logarithm_table[7041] = 14'b0000101_1100100;
		logarithm_table[7042] = 14'b0000101_1100100;
		logarithm_table[7043] = 14'b0000101_1100100;
		logarithm_table[7044] = 14'b0000101_1100100;
		logarithm_table[7045] = 14'b0000101_1100100;
		logarithm_table[7046] = 14'b0000101_1100100;
		logarithm_table[7047] = 14'b0000101_1100100;
		logarithm_table[7048] = 14'b0000101_1100100;
		logarithm_table[7049] = 14'b0000101_1100100;
		logarithm_table[7050] = 14'b0000101_1100100;
		logarithm_table[7051] = 14'b0000101_1100100;
		logarithm_table[7052] = 14'b0000101_1100100;
		logarithm_table[7053] = 14'b0000101_1100100;
		logarithm_table[7054] = 14'b0000101_1100100;
		logarithm_table[7055] = 14'b0000101_1100100;
		logarithm_table[7056] = 14'b0000101_1100100;
		logarithm_table[7057] = 14'b0000101_1100100;
		logarithm_table[7058] = 14'b0000101_1100100;
		logarithm_table[7059] = 14'b0000101_1100101;
		logarithm_table[7060] = 14'b0000101_1100101;
		logarithm_table[7061] = 14'b0000101_1100101;
		logarithm_table[7062] = 14'b0000101_1100101;
		logarithm_table[7063] = 14'b0000101_1100101;
		logarithm_table[7064] = 14'b0000101_1100101;
		logarithm_table[7065] = 14'b0000101_1100101;
		logarithm_table[7066] = 14'b0000101_1100101;
		logarithm_table[7067] = 14'b0000101_1100101;
		logarithm_table[7068] = 14'b0000101_1100101;
		logarithm_table[7069] = 14'b0000101_1100101;
		logarithm_table[7070] = 14'b0000101_1100101;
		logarithm_table[7071] = 14'b0000101_1100101;
		logarithm_table[7072] = 14'b0000101_1100101;
		logarithm_table[7073] = 14'b0000101_1100101;
		logarithm_table[7074] = 14'b0000101_1100101;
		logarithm_table[7075] = 14'b0000101_1100101;
		logarithm_table[7076] = 14'b0000101_1100101;
		logarithm_table[7077] = 14'b0000101_1100101;
		logarithm_table[7078] = 14'b0000101_1100101;
		logarithm_table[7079] = 14'b0000101_1100101;
		logarithm_table[7080] = 14'b0000101_1100101;
		logarithm_table[7081] = 14'b0000101_1100101;
		logarithm_table[7082] = 14'b0000101_1100101;
		logarithm_table[7083] = 14'b0000101_1100101;
		logarithm_table[7084] = 14'b0000101_1100101;
		logarithm_table[7085] = 14'b0000101_1100101;
		logarithm_table[7086] = 14'b0000101_1100101;
		logarithm_table[7087] = 14'b0000101_1100101;
		logarithm_table[7088] = 14'b0000101_1100101;
		logarithm_table[7089] = 14'b0000101_1100101;
		logarithm_table[7090] = 14'b0000101_1100101;
		logarithm_table[7091] = 14'b0000101_1100101;
		logarithm_table[7092] = 14'b0000101_1100101;
		logarithm_table[7093] = 14'b0000101_1100101;
		logarithm_table[7094] = 14'b0000101_1100101;
		logarithm_table[7095] = 14'b0000101_1100101;
		logarithm_table[7096] = 14'b0000101_1100101;
		logarithm_table[7097] = 14'b0000101_1100110;
		logarithm_table[7098] = 14'b0000101_1100110;
		logarithm_table[7099] = 14'b0000101_1100110;
		logarithm_table[7100] = 14'b0000101_1100110;
		logarithm_table[7101] = 14'b0000101_1100110;
		logarithm_table[7102] = 14'b0000101_1100110;
		logarithm_table[7103] = 14'b0000101_1100110;
		logarithm_table[7104] = 14'b0000101_1100110;
		logarithm_table[7105] = 14'b0000101_1100110;
		logarithm_table[7106] = 14'b0000101_1100110;
		logarithm_table[7107] = 14'b0000101_1100110;
		logarithm_table[7108] = 14'b0000101_1100110;
		logarithm_table[7109] = 14'b0000101_1100110;
		logarithm_table[7110] = 14'b0000101_1100110;
		logarithm_table[7111] = 14'b0000101_1100110;
		logarithm_table[7112] = 14'b0000101_1100110;
		logarithm_table[7113] = 14'b0000101_1100110;
		logarithm_table[7114] = 14'b0000101_1100110;
		logarithm_table[7115] = 14'b0000101_1100110;
		logarithm_table[7116] = 14'b0000101_1100110;
		logarithm_table[7117] = 14'b0000101_1100110;
		logarithm_table[7118] = 14'b0000101_1100110;
		logarithm_table[7119] = 14'b0000101_1100110;
		logarithm_table[7120] = 14'b0000101_1100110;
		logarithm_table[7121] = 14'b0000101_1100110;
		logarithm_table[7122] = 14'b0000101_1100110;
		logarithm_table[7123] = 14'b0000101_1100110;
		logarithm_table[7124] = 14'b0000101_1100110;
		logarithm_table[7125] = 14'b0000101_1100110;
		logarithm_table[7126] = 14'b0000101_1100110;
		logarithm_table[7127] = 14'b0000101_1100110;
		logarithm_table[7128] = 14'b0000101_1100110;
		logarithm_table[7129] = 14'b0000101_1100110;
		logarithm_table[7130] = 14'b0000101_1100110;
		logarithm_table[7131] = 14'b0000101_1100110;
		logarithm_table[7132] = 14'b0000101_1100110;
		logarithm_table[7133] = 14'b0000101_1100110;
		logarithm_table[7134] = 14'b0000101_1100110;
		logarithm_table[7135] = 14'b0000101_1100110;
		logarithm_table[7136] = 14'b0000101_1100111;
		logarithm_table[7137] = 14'b0000101_1100111;
		logarithm_table[7138] = 14'b0000101_1100111;
		logarithm_table[7139] = 14'b0000101_1100111;
		logarithm_table[7140] = 14'b0000101_1100111;
		logarithm_table[7141] = 14'b0000101_1100111;
		logarithm_table[7142] = 14'b0000101_1100111;
		logarithm_table[7143] = 14'b0000101_1100111;
		logarithm_table[7144] = 14'b0000101_1100111;
		logarithm_table[7145] = 14'b0000101_1100111;
		logarithm_table[7146] = 14'b0000101_1100111;
		logarithm_table[7147] = 14'b0000101_1100111;
		logarithm_table[7148] = 14'b0000101_1100111;
		logarithm_table[7149] = 14'b0000101_1100111;
		logarithm_table[7150] = 14'b0000101_1100111;
		logarithm_table[7151] = 14'b0000101_1100111;
		logarithm_table[7152] = 14'b0000101_1100111;
		logarithm_table[7153] = 14'b0000101_1100111;
		logarithm_table[7154] = 14'b0000101_1100111;
		logarithm_table[7155] = 14'b0000101_1100111;
		logarithm_table[7156] = 14'b0000101_1100111;
		logarithm_table[7157] = 14'b0000101_1100111;
		logarithm_table[7158] = 14'b0000101_1100111;
		logarithm_table[7159] = 14'b0000101_1100111;
		logarithm_table[7160] = 14'b0000101_1100111;
		logarithm_table[7161] = 14'b0000101_1100111;
		logarithm_table[7162] = 14'b0000101_1100111;
		logarithm_table[7163] = 14'b0000101_1100111;
		logarithm_table[7164] = 14'b0000101_1100111;
		logarithm_table[7165] = 14'b0000101_1100111;
		logarithm_table[7166] = 14'b0000101_1100111;
		logarithm_table[7167] = 14'b0000101_1100111;
		logarithm_table[7168] = 14'b0000101_1100111;
		logarithm_table[7169] = 14'b0000101_1100111;
		logarithm_table[7170] = 14'b0000101_1100111;
		logarithm_table[7171] = 14'b0000101_1100111;
		logarithm_table[7172] = 14'b0000101_1100111;
		logarithm_table[7173] = 14'b0000101_1100111;
		logarithm_table[7174] = 14'b0000101_1100111;
		logarithm_table[7175] = 14'b0000101_1101000;
		logarithm_table[7176] = 14'b0000101_1101000;
		logarithm_table[7177] = 14'b0000101_1101000;
		logarithm_table[7178] = 14'b0000101_1101000;
		logarithm_table[7179] = 14'b0000101_1101000;
		logarithm_table[7180] = 14'b0000101_1101000;
		logarithm_table[7181] = 14'b0000101_1101000;
		logarithm_table[7182] = 14'b0000101_1101000;
		logarithm_table[7183] = 14'b0000101_1101000;
		logarithm_table[7184] = 14'b0000101_1101000;
		logarithm_table[7185] = 14'b0000101_1101000;
		logarithm_table[7186] = 14'b0000101_1101000;
		logarithm_table[7187] = 14'b0000101_1101000;
		logarithm_table[7188] = 14'b0000101_1101000;
		logarithm_table[7189] = 14'b0000101_1101000;
		logarithm_table[7190] = 14'b0000101_1101000;
		logarithm_table[7191] = 14'b0000101_1101000;
		logarithm_table[7192] = 14'b0000101_1101000;
		logarithm_table[7193] = 14'b0000101_1101000;
		logarithm_table[7194] = 14'b0000101_1101000;
		logarithm_table[7195] = 14'b0000101_1101000;
		logarithm_table[7196] = 14'b0000101_1101000;
		logarithm_table[7197] = 14'b0000101_1101000;
		logarithm_table[7198] = 14'b0000101_1101000;
		logarithm_table[7199] = 14'b0000101_1101000;
		logarithm_table[7200] = 14'b0000101_1101000;
		logarithm_table[7201] = 14'b0000101_1101000;
		logarithm_table[7202] = 14'b0000101_1101000;
		logarithm_table[7203] = 14'b0000101_1101000;
		logarithm_table[7204] = 14'b0000101_1101000;
		logarithm_table[7205] = 14'b0000101_1101000;
		logarithm_table[7206] = 14'b0000101_1101000;
		logarithm_table[7207] = 14'b0000101_1101000;
		logarithm_table[7208] = 14'b0000101_1101000;
		logarithm_table[7209] = 14'b0000101_1101000;
		logarithm_table[7210] = 14'b0000101_1101000;
		logarithm_table[7211] = 14'b0000101_1101000;
		logarithm_table[7212] = 14'b0000101_1101000;
		logarithm_table[7213] = 14'b0000101_1101000;
		logarithm_table[7214] = 14'b0000101_1101001;
		logarithm_table[7215] = 14'b0000101_1101001;
		logarithm_table[7216] = 14'b0000101_1101001;
		logarithm_table[7217] = 14'b0000101_1101001;
		logarithm_table[7218] = 14'b0000101_1101001;
		logarithm_table[7219] = 14'b0000101_1101001;
		logarithm_table[7220] = 14'b0000101_1101001;
		logarithm_table[7221] = 14'b0000101_1101001;
		logarithm_table[7222] = 14'b0000101_1101001;
		logarithm_table[7223] = 14'b0000101_1101001;
		logarithm_table[7224] = 14'b0000101_1101001;
		logarithm_table[7225] = 14'b0000101_1101001;
		logarithm_table[7226] = 14'b0000101_1101001;
		logarithm_table[7227] = 14'b0000101_1101001;
		logarithm_table[7228] = 14'b0000101_1101001;
		logarithm_table[7229] = 14'b0000101_1101001;
		logarithm_table[7230] = 14'b0000101_1101001;
		logarithm_table[7231] = 14'b0000101_1101001;
		logarithm_table[7232] = 14'b0000101_1101001;
		logarithm_table[7233] = 14'b0000101_1101001;
		logarithm_table[7234] = 14'b0000101_1101001;
		logarithm_table[7235] = 14'b0000101_1101001;
		logarithm_table[7236] = 14'b0000101_1101001;
		logarithm_table[7237] = 14'b0000101_1101001;
		logarithm_table[7238] = 14'b0000101_1101001;
		logarithm_table[7239] = 14'b0000101_1101001;
		logarithm_table[7240] = 14'b0000101_1101001;
		logarithm_table[7241] = 14'b0000101_1101001;
		logarithm_table[7242] = 14'b0000101_1101001;
		logarithm_table[7243] = 14'b0000101_1101001;
		logarithm_table[7244] = 14'b0000101_1101001;
		logarithm_table[7245] = 14'b0000101_1101001;
		logarithm_table[7246] = 14'b0000101_1101001;
		logarithm_table[7247] = 14'b0000101_1101001;
		logarithm_table[7248] = 14'b0000101_1101001;
		logarithm_table[7249] = 14'b0000101_1101001;
		logarithm_table[7250] = 14'b0000101_1101001;
		logarithm_table[7251] = 14'b0000101_1101001;
		logarithm_table[7252] = 14'b0000101_1101001;
		logarithm_table[7253] = 14'b0000101_1101010;
		logarithm_table[7254] = 14'b0000101_1101010;
		logarithm_table[7255] = 14'b0000101_1101010;
		logarithm_table[7256] = 14'b0000101_1101010;
		logarithm_table[7257] = 14'b0000101_1101010;
		logarithm_table[7258] = 14'b0000101_1101010;
		logarithm_table[7259] = 14'b0000101_1101010;
		logarithm_table[7260] = 14'b0000101_1101010;
		logarithm_table[7261] = 14'b0000101_1101010;
		logarithm_table[7262] = 14'b0000101_1101010;
		logarithm_table[7263] = 14'b0000101_1101010;
		logarithm_table[7264] = 14'b0000101_1101010;
		logarithm_table[7265] = 14'b0000101_1101010;
		logarithm_table[7266] = 14'b0000101_1101010;
		logarithm_table[7267] = 14'b0000101_1101010;
		logarithm_table[7268] = 14'b0000101_1101010;
		logarithm_table[7269] = 14'b0000101_1101010;
		logarithm_table[7270] = 14'b0000101_1101010;
		logarithm_table[7271] = 14'b0000101_1101010;
		logarithm_table[7272] = 14'b0000101_1101010;
		logarithm_table[7273] = 14'b0000101_1101010;
		logarithm_table[7274] = 14'b0000101_1101010;
		logarithm_table[7275] = 14'b0000101_1101010;
		logarithm_table[7276] = 14'b0000101_1101010;
		logarithm_table[7277] = 14'b0000101_1101010;
		logarithm_table[7278] = 14'b0000101_1101010;
		logarithm_table[7279] = 14'b0000101_1101010;
		logarithm_table[7280] = 14'b0000101_1101010;
		logarithm_table[7281] = 14'b0000101_1101010;
		logarithm_table[7282] = 14'b0000101_1101010;
		logarithm_table[7283] = 14'b0000101_1101010;
		logarithm_table[7284] = 14'b0000101_1101010;
		logarithm_table[7285] = 14'b0000101_1101010;
		logarithm_table[7286] = 14'b0000101_1101010;
		logarithm_table[7287] = 14'b0000101_1101010;
		logarithm_table[7288] = 14'b0000101_1101010;
		logarithm_table[7289] = 14'b0000101_1101010;
		logarithm_table[7290] = 14'b0000101_1101010;
		logarithm_table[7291] = 14'b0000101_1101010;
		logarithm_table[7292] = 14'b0000101_1101011;
		logarithm_table[7293] = 14'b0000101_1101011;
		logarithm_table[7294] = 14'b0000101_1101011;
		logarithm_table[7295] = 14'b0000101_1101011;
		logarithm_table[7296] = 14'b0000101_1101011;
		logarithm_table[7297] = 14'b0000101_1101011;
		logarithm_table[7298] = 14'b0000101_1101011;
		logarithm_table[7299] = 14'b0000101_1101011;
		logarithm_table[7300] = 14'b0000101_1101011;
		logarithm_table[7301] = 14'b0000101_1101011;
		logarithm_table[7302] = 14'b0000101_1101011;
		logarithm_table[7303] = 14'b0000101_1101011;
		logarithm_table[7304] = 14'b0000101_1101011;
		logarithm_table[7305] = 14'b0000101_1101011;
		logarithm_table[7306] = 14'b0000101_1101011;
		logarithm_table[7307] = 14'b0000101_1101011;
		logarithm_table[7308] = 14'b0000101_1101011;
		logarithm_table[7309] = 14'b0000101_1101011;
		logarithm_table[7310] = 14'b0000101_1101011;
		logarithm_table[7311] = 14'b0000101_1101011;
		logarithm_table[7312] = 14'b0000101_1101011;
		logarithm_table[7313] = 14'b0000101_1101011;
		logarithm_table[7314] = 14'b0000101_1101011;
		logarithm_table[7315] = 14'b0000101_1101011;
		logarithm_table[7316] = 14'b0000101_1101011;
		logarithm_table[7317] = 14'b0000101_1101011;
		logarithm_table[7318] = 14'b0000101_1101011;
		logarithm_table[7319] = 14'b0000101_1101011;
		logarithm_table[7320] = 14'b0000101_1101011;
		logarithm_table[7321] = 14'b0000101_1101011;
		logarithm_table[7322] = 14'b0000101_1101011;
		logarithm_table[7323] = 14'b0000101_1101011;
		logarithm_table[7324] = 14'b0000101_1101011;
		logarithm_table[7325] = 14'b0000101_1101011;
		logarithm_table[7326] = 14'b0000101_1101011;
		logarithm_table[7327] = 14'b0000101_1101011;
		logarithm_table[7328] = 14'b0000101_1101011;
		logarithm_table[7329] = 14'b0000101_1101011;
		logarithm_table[7330] = 14'b0000101_1101011;
		logarithm_table[7331] = 14'b0000101_1101011;
		logarithm_table[7332] = 14'b0000101_1101100;
		logarithm_table[7333] = 14'b0000101_1101100;
		logarithm_table[7334] = 14'b0000101_1101100;
		logarithm_table[7335] = 14'b0000101_1101100;
		logarithm_table[7336] = 14'b0000101_1101100;
		logarithm_table[7337] = 14'b0000101_1101100;
		logarithm_table[7338] = 14'b0000101_1101100;
		logarithm_table[7339] = 14'b0000101_1101100;
		logarithm_table[7340] = 14'b0000101_1101100;
		logarithm_table[7341] = 14'b0000101_1101100;
		logarithm_table[7342] = 14'b0000101_1101100;
		logarithm_table[7343] = 14'b0000101_1101100;
		logarithm_table[7344] = 14'b0000101_1101100;
		logarithm_table[7345] = 14'b0000101_1101100;
		logarithm_table[7346] = 14'b0000101_1101100;
		logarithm_table[7347] = 14'b0000101_1101100;
		logarithm_table[7348] = 14'b0000101_1101100;
		logarithm_table[7349] = 14'b0000101_1101100;
		logarithm_table[7350] = 14'b0000101_1101100;
		logarithm_table[7351] = 14'b0000101_1101100;
		logarithm_table[7352] = 14'b0000101_1101100;
		logarithm_table[7353] = 14'b0000101_1101100;
		logarithm_table[7354] = 14'b0000101_1101100;
		logarithm_table[7355] = 14'b0000101_1101100;
		logarithm_table[7356] = 14'b0000101_1101100;
		logarithm_table[7357] = 14'b0000101_1101100;
		logarithm_table[7358] = 14'b0000101_1101100;
		logarithm_table[7359] = 14'b0000101_1101100;
		logarithm_table[7360] = 14'b0000101_1101100;
		logarithm_table[7361] = 14'b0000101_1101100;
		logarithm_table[7362] = 14'b0000101_1101100;
		logarithm_table[7363] = 14'b0000101_1101100;
		logarithm_table[7364] = 14'b0000101_1101100;
		logarithm_table[7365] = 14'b0000101_1101100;
		logarithm_table[7366] = 14'b0000101_1101100;
		logarithm_table[7367] = 14'b0000101_1101100;
		logarithm_table[7368] = 14'b0000101_1101100;
		logarithm_table[7369] = 14'b0000101_1101100;
		logarithm_table[7370] = 14'b0000101_1101100;
		logarithm_table[7371] = 14'b0000101_1101100;
		logarithm_table[7372] = 14'b0000101_1101101;
		logarithm_table[7373] = 14'b0000101_1101101;
		logarithm_table[7374] = 14'b0000101_1101101;
		logarithm_table[7375] = 14'b0000101_1101101;
		logarithm_table[7376] = 14'b0000101_1101101;
		logarithm_table[7377] = 14'b0000101_1101101;
		logarithm_table[7378] = 14'b0000101_1101101;
		logarithm_table[7379] = 14'b0000101_1101101;
		logarithm_table[7380] = 14'b0000101_1101101;
		logarithm_table[7381] = 14'b0000101_1101101;
		logarithm_table[7382] = 14'b0000101_1101101;
		logarithm_table[7383] = 14'b0000101_1101101;
		logarithm_table[7384] = 14'b0000101_1101101;
		logarithm_table[7385] = 14'b0000101_1101101;
		logarithm_table[7386] = 14'b0000101_1101101;
		logarithm_table[7387] = 14'b0000101_1101101;
		logarithm_table[7388] = 14'b0000101_1101101;
		logarithm_table[7389] = 14'b0000101_1101101;
		logarithm_table[7390] = 14'b0000101_1101101;
		logarithm_table[7391] = 14'b0000101_1101101;
		logarithm_table[7392] = 14'b0000101_1101101;
		logarithm_table[7393] = 14'b0000101_1101101;
		logarithm_table[7394] = 14'b0000101_1101101;
		logarithm_table[7395] = 14'b0000101_1101101;
		logarithm_table[7396] = 14'b0000101_1101101;
		logarithm_table[7397] = 14'b0000101_1101101;
		logarithm_table[7398] = 14'b0000101_1101101;
		logarithm_table[7399] = 14'b0000101_1101101;
		logarithm_table[7400] = 14'b0000101_1101101;
		logarithm_table[7401] = 14'b0000101_1101101;
		logarithm_table[7402] = 14'b0000101_1101101;
		logarithm_table[7403] = 14'b0000101_1101101;
		logarithm_table[7404] = 14'b0000101_1101101;
		logarithm_table[7405] = 14'b0000101_1101101;
		logarithm_table[7406] = 14'b0000101_1101101;
		logarithm_table[7407] = 14'b0000101_1101101;
		logarithm_table[7408] = 14'b0000101_1101101;
		logarithm_table[7409] = 14'b0000101_1101101;
		logarithm_table[7410] = 14'b0000101_1101101;
		logarithm_table[7411] = 14'b0000101_1101101;
		logarithm_table[7412] = 14'b0000101_1101110;
		logarithm_table[7413] = 14'b0000101_1101110;
		logarithm_table[7414] = 14'b0000101_1101110;
		logarithm_table[7415] = 14'b0000101_1101110;
		logarithm_table[7416] = 14'b0000101_1101110;
		logarithm_table[7417] = 14'b0000101_1101110;
		logarithm_table[7418] = 14'b0000101_1101110;
		logarithm_table[7419] = 14'b0000101_1101110;
		logarithm_table[7420] = 14'b0000101_1101110;
		logarithm_table[7421] = 14'b0000101_1101110;
		logarithm_table[7422] = 14'b0000101_1101110;
		logarithm_table[7423] = 14'b0000101_1101110;
		logarithm_table[7424] = 14'b0000101_1101110;
		logarithm_table[7425] = 14'b0000101_1101110;
		logarithm_table[7426] = 14'b0000101_1101110;
		logarithm_table[7427] = 14'b0000101_1101110;
		logarithm_table[7428] = 14'b0000101_1101110;
		logarithm_table[7429] = 14'b0000101_1101110;
		logarithm_table[7430] = 14'b0000101_1101110;
		logarithm_table[7431] = 14'b0000101_1101110;
		logarithm_table[7432] = 14'b0000101_1101110;
		logarithm_table[7433] = 14'b0000101_1101110;
		logarithm_table[7434] = 14'b0000101_1101110;
		logarithm_table[7435] = 14'b0000101_1101110;
		logarithm_table[7436] = 14'b0000101_1101110;
		logarithm_table[7437] = 14'b0000101_1101110;
		logarithm_table[7438] = 14'b0000101_1101110;
		logarithm_table[7439] = 14'b0000101_1101110;
		logarithm_table[7440] = 14'b0000101_1101110;
		logarithm_table[7441] = 14'b0000101_1101110;
		logarithm_table[7442] = 14'b0000101_1101110;
		logarithm_table[7443] = 14'b0000101_1101110;
		logarithm_table[7444] = 14'b0000101_1101110;
		logarithm_table[7445] = 14'b0000101_1101110;
		logarithm_table[7446] = 14'b0000101_1101110;
		logarithm_table[7447] = 14'b0000101_1101110;
		logarithm_table[7448] = 14'b0000101_1101110;
		logarithm_table[7449] = 14'b0000101_1101110;
		logarithm_table[7450] = 14'b0000101_1101110;
		logarithm_table[7451] = 14'b0000101_1101110;
		logarithm_table[7452] = 14'b0000101_1101111;
		logarithm_table[7453] = 14'b0000101_1101111;
		logarithm_table[7454] = 14'b0000101_1101111;
		logarithm_table[7455] = 14'b0000101_1101111;
		logarithm_table[7456] = 14'b0000101_1101111;
		logarithm_table[7457] = 14'b0000101_1101111;
		logarithm_table[7458] = 14'b0000101_1101111;
		logarithm_table[7459] = 14'b0000101_1101111;
		logarithm_table[7460] = 14'b0000101_1101111;
		logarithm_table[7461] = 14'b0000101_1101111;
		logarithm_table[7462] = 14'b0000101_1101111;
		logarithm_table[7463] = 14'b0000101_1101111;
		logarithm_table[7464] = 14'b0000101_1101111;
		logarithm_table[7465] = 14'b0000101_1101111;
		logarithm_table[7466] = 14'b0000101_1101111;
		logarithm_table[7467] = 14'b0000101_1101111;
		logarithm_table[7468] = 14'b0000101_1101111;
		logarithm_table[7469] = 14'b0000101_1101111;
		logarithm_table[7470] = 14'b0000101_1101111;
		logarithm_table[7471] = 14'b0000101_1101111;
		logarithm_table[7472] = 14'b0000101_1101111;
		logarithm_table[7473] = 14'b0000101_1101111;
		logarithm_table[7474] = 14'b0000101_1101111;
		logarithm_table[7475] = 14'b0000101_1101111;
		logarithm_table[7476] = 14'b0000101_1101111;
		logarithm_table[7477] = 14'b0000101_1101111;
		logarithm_table[7478] = 14'b0000101_1101111;
		logarithm_table[7479] = 14'b0000101_1101111;
		logarithm_table[7480] = 14'b0000101_1101111;
		logarithm_table[7481] = 14'b0000101_1101111;
		logarithm_table[7482] = 14'b0000101_1101111;
		logarithm_table[7483] = 14'b0000101_1101111;
		logarithm_table[7484] = 14'b0000101_1101111;
		logarithm_table[7485] = 14'b0000101_1101111;
		logarithm_table[7486] = 14'b0000101_1101111;
		logarithm_table[7487] = 14'b0000101_1101111;
		logarithm_table[7488] = 14'b0000101_1101111;
		logarithm_table[7489] = 14'b0000101_1101111;
		logarithm_table[7490] = 14'b0000101_1101111;
		logarithm_table[7491] = 14'b0000101_1101111;
		logarithm_table[7492] = 14'b0000101_1110000;
		logarithm_table[7493] = 14'b0000101_1110000;
		logarithm_table[7494] = 14'b0000101_1110000;
		logarithm_table[7495] = 14'b0000101_1110000;
		logarithm_table[7496] = 14'b0000101_1110000;
		logarithm_table[7497] = 14'b0000101_1110000;
		logarithm_table[7498] = 14'b0000101_1110000;
		logarithm_table[7499] = 14'b0000101_1110000;
		logarithm_table[7500] = 14'b0000101_1110000;
		logarithm_table[7501] = 14'b0000101_1110000;
		logarithm_table[7502] = 14'b0000101_1110000;
		logarithm_table[7503] = 14'b0000101_1110000;
		logarithm_table[7504] = 14'b0000101_1110000;
		logarithm_table[7505] = 14'b0000101_1110000;
		logarithm_table[7506] = 14'b0000101_1110000;
		logarithm_table[7507] = 14'b0000101_1110000;
		logarithm_table[7508] = 14'b0000101_1110000;
		logarithm_table[7509] = 14'b0000101_1110000;
		logarithm_table[7510] = 14'b0000101_1110000;
		logarithm_table[7511] = 14'b0000101_1110000;
		logarithm_table[7512] = 14'b0000101_1110000;
		logarithm_table[7513] = 14'b0000101_1110000;
		logarithm_table[7514] = 14'b0000101_1110000;
		logarithm_table[7515] = 14'b0000101_1110000;
		logarithm_table[7516] = 14'b0000101_1110000;
		logarithm_table[7517] = 14'b0000101_1110000;
		logarithm_table[7518] = 14'b0000101_1110000;
		logarithm_table[7519] = 14'b0000101_1110000;
		logarithm_table[7520] = 14'b0000101_1110000;
		logarithm_table[7521] = 14'b0000101_1110000;
		logarithm_table[7522] = 14'b0000101_1110000;
		logarithm_table[7523] = 14'b0000101_1110000;
		logarithm_table[7524] = 14'b0000101_1110000;
		logarithm_table[7525] = 14'b0000101_1110000;
		logarithm_table[7526] = 14'b0000101_1110000;
		logarithm_table[7527] = 14'b0000101_1110000;
		logarithm_table[7528] = 14'b0000101_1110000;
		logarithm_table[7529] = 14'b0000101_1110000;
		logarithm_table[7530] = 14'b0000101_1110000;
		logarithm_table[7531] = 14'b0000101_1110000;
		logarithm_table[7532] = 14'b0000101_1110000;
		logarithm_table[7533] = 14'b0000101_1110001;
		logarithm_table[7534] = 14'b0000101_1110001;
		logarithm_table[7535] = 14'b0000101_1110001;
		logarithm_table[7536] = 14'b0000101_1110001;
		logarithm_table[7537] = 14'b0000101_1110001;
		logarithm_table[7538] = 14'b0000101_1110001;
		logarithm_table[7539] = 14'b0000101_1110001;
		logarithm_table[7540] = 14'b0000101_1110001;
		logarithm_table[7541] = 14'b0000101_1110001;
		logarithm_table[7542] = 14'b0000101_1110001;
		logarithm_table[7543] = 14'b0000101_1110001;
		logarithm_table[7544] = 14'b0000101_1110001;
		logarithm_table[7545] = 14'b0000101_1110001;
		logarithm_table[7546] = 14'b0000101_1110001;
		logarithm_table[7547] = 14'b0000101_1110001;
		logarithm_table[7548] = 14'b0000101_1110001;
		logarithm_table[7549] = 14'b0000101_1110001;
		logarithm_table[7550] = 14'b0000101_1110001;
		logarithm_table[7551] = 14'b0000101_1110001;
		logarithm_table[7552] = 14'b0000101_1110001;
		logarithm_table[7553] = 14'b0000101_1110001;
		logarithm_table[7554] = 14'b0000101_1110001;
		logarithm_table[7555] = 14'b0000101_1110001;
		logarithm_table[7556] = 14'b0000101_1110001;
		logarithm_table[7557] = 14'b0000101_1110001;
		logarithm_table[7558] = 14'b0000101_1110001;
		logarithm_table[7559] = 14'b0000101_1110001;
		logarithm_table[7560] = 14'b0000101_1110001;
		logarithm_table[7561] = 14'b0000101_1110001;
		logarithm_table[7562] = 14'b0000101_1110001;
		logarithm_table[7563] = 14'b0000101_1110001;
		logarithm_table[7564] = 14'b0000101_1110001;
		logarithm_table[7565] = 14'b0000101_1110001;
		logarithm_table[7566] = 14'b0000101_1110001;
		logarithm_table[7567] = 14'b0000101_1110001;
		logarithm_table[7568] = 14'b0000101_1110001;
		logarithm_table[7569] = 14'b0000101_1110001;
		logarithm_table[7570] = 14'b0000101_1110001;
		logarithm_table[7571] = 14'b0000101_1110001;
		logarithm_table[7572] = 14'b0000101_1110001;
		logarithm_table[7573] = 14'b0000101_1110001;
		logarithm_table[7574] = 14'b0000101_1110010;
		logarithm_table[7575] = 14'b0000101_1110010;
		logarithm_table[7576] = 14'b0000101_1110010;
		logarithm_table[7577] = 14'b0000101_1110010;
		logarithm_table[7578] = 14'b0000101_1110010;
		logarithm_table[7579] = 14'b0000101_1110010;
		logarithm_table[7580] = 14'b0000101_1110010;
		logarithm_table[7581] = 14'b0000101_1110010;
		logarithm_table[7582] = 14'b0000101_1110010;
		logarithm_table[7583] = 14'b0000101_1110010;
		logarithm_table[7584] = 14'b0000101_1110010;
		logarithm_table[7585] = 14'b0000101_1110010;
		logarithm_table[7586] = 14'b0000101_1110010;
		logarithm_table[7587] = 14'b0000101_1110010;
		logarithm_table[7588] = 14'b0000101_1110010;
		logarithm_table[7589] = 14'b0000101_1110010;
		logarithm_table[7590] = 14'b0000101_1110010;
		logarithm_table[7591] = 14'b0000101_1110010;
		logarithm_table[7592] = 14'b0000101_1110010;
		logarithm_table[7593] = 14'b0000101_1110010;
		logarithm_table[7594] = 14'b0000101_1110010;
		logarithm_table[7595] = 14'b0000101_1110010;
		logarithm_table[7596] = 14'b0000101_1110010;
		logarithm_table[7597] = 14'b0000101_1110010;
		logarithm_table[7598] = 14'b0000101_1110010;
		logarithm_table[7599] = 14'b0000101_1110010;
		logarithm_table[7600] = 14'b0000101_1110010;
		logarithm_table[7601] = 14'b0000101_1110010;
		logarithm_table[7602] = 14'b0000101_1110010;
		logarithm_table[7603] = 14'b0000101_1110010;
		logarithm_table[7604] = 14'b0000101_1110010;
		logarithm_table[7605] = 14'b0000101_1110010;
		logarithm_table[7606] = 14'b0000101_1110010;
		logarithm_table[7607] = 14'b0000101_1110010;
		logarithm_table[7608] = 14'b0000101_1110010;
		logarithm_table[7609] = 14'b0000101_1110010;
		logarithm_table[7610] = 14'b0000101_1110010;
		logarithm_table[7611] = 14'b0000101_1110010;
		logarithm_table[7612] = 14'b0000101_1110010;
		logarithm_table[7613] = 14'b0000101_1110010;
		logarithm_table[7614] = 14'b0000101_1110010;
		logarithm_table[7615] = 14'b0000101_1110011;
		logarithm_table[7616] = 14'b0000101_1110011;
		logarithm_table[7617] = 14'b0000101_1110011;
		logarithm_table[7618] = 14'b0000101_1110011;
		logarithm_table[7619] = 14'b0000101_1110011;
		logarithm_table[7620] = 14'b0000101_1110011;
		logarithm_table[7621] = 14'b0000101_1110011;
		logarithm_table[7622] = 14'b0000101_1110011;
		logarithm_table[7623] = 14'b0000101_1110011;
		logarithm_table[7624] = 14'b0000101_1110011;
		logarithm_table[7625] = 14'b0000101_1110011;
		logarithm_table[7626] = 14'b0000101_1110011;
		logarithm_table[7627] = 14'b0000101_1110011;
		logarithm_table[7628] = 14'b0000101_1110011;
		logarithm_table[7629] = 14'b0000101_1110011;
		logarithm_table[7630] = 14'b0000101_1110011;
		logarithm_table[7631] = 14'b0000101_1110011;
		logarithm_table[7632] = 14'b0000101_1110011;
		logarithm_table[7633] = 14'b0000101_1110011;
		logarithm_table[7634] = 14'b0000101_1110011;
		logarithm_table[7635] = 14'b0000101_1110011;
		logarithm_table[7636] = 14'b0000101_1110011;
		logarithm_table[7637] = 14'b0000101_1110011;
		logarithm_table[7638] = 14'b0000101_1110011;
		logarithm_table[7639] = 14'b0000101_1110011;
		logarithm_table[7640] = 14'b0000101_1110011;
		logarithm_table[7641] = 14'b0000101_1110011;
		logarithm_table[7642] = 14'b0000101_1110011;
		logarithm_table[7643] = 14'b0000101_1110011;
		logarithm_table[7644] = 14'b0000101_1110011;
		logarithm_table[7645] = 14'b0000101_1110011;
		logarithm_table[7646] = 14'b0000101_1110011;
		logarithm_table[7647] = 14'b0000101_1110011;
		logarithm_table[7648] = 14'b0000101_1110011;
		logarithm_table[7649] = 14'b0000101_1110011;
		logarithm_table[7650] = 14'b0000101_1110011;
		logarithm_table[7651] = 14'b0000101_1110011;
		logarithm_table[7652] = 14'b0000101_1110011;
		logarithm_table[7653] = 14'b0000101_1110011;
		logarithm_table[7654] = 14'b0000101_1110011;
		logarithm_table[7655] = 14'b0000101_1110011;
		logarithm_table[7656] = 14'b0000101_1110100;
		logarithm_table[7657] = 14'b0000101_1110100;
		logarithm_table[7658] = 14'b0000101_1110100;
		logarithm_table[7659] = 14'b0000101_1110100;
		logarithm_table[7660] = 14'b0000101_1110100;
		logarithm_table[7661] = 14'b0000101_1110100;
		logarithm_table[7662] = 14'b0000101_1110100;
		logarithm_table[7663] = 14'b0000101_1110100;
		logarithm_table[7664] = 14'b0000101_1110100;
		logarithm_table[7665] = 14'b0000101_1110100;
		logarithm_table[7666] = 14'b0000101_1110100;
		logarithm_table[7667] = 14'b0000101_1110100;
		logarithm_table[7668] = 14'b0000101_1110100;
		logarithm_table[7669] = 14'b0000101_1110100;
		logarithm_table[7670] = 14'b0000101_1110100;
		logarithm_table[7671] = 14'b0000101_1110100;
		logarithm_table[7672] = 14'b0000101_1110100;
		logarithm_table[7673] = 14'b0000101_1110100;
		logarithm_table[7674] = 14'b0000101_1110100;
		logarithm_table[7675] = 14'b0000101_1110100;
		logarithm_table[7676] = 14'b0000101_1110100;
		logarithm_table[7677] = 14'b0000101_1110100;
		logarithm_table[7678] = 14'b0000101_1110100;
		logarithm_table[7679] = 14'b0000101_1110100;
		logarithm_table[7680] = 14'b0000101_1110100;
		logarithm_table[7681] = 14'b0000101_1110100;
		logarithm_table[7682] = 14'b0000101_1110100;
		logarithm_table[7683] = 14'b0000101_1110100;
		logarithm_table[7684] = 14'b0000101_1110100;
		logarithm_table[7685] = 14'b0000101_1110100;
		logarithm_table[7686] = 14'b0000101_1110100;
		logarithm_table[7687] = 14'b0000101_1110100;
		logarithm_table[7688] = 14'b0000101_1110100;
		logarithm_table[7689] = 14'b0000101_1110100;
		logarithm_table[7690] = 14'b0000101_1110100;
		logarithm_table[7691] = 14'b0000101_1110100;
		logarithm_table[7692] = 14'b0000101_1110100;
		logarithm_table[7693] = 14'b0000101_1110100;
		logarithm_table[7694] = 14'b0000101_1110100;
		logarithm_table[7695] = 14'b0000101_1110100;
		logarithm_table[7696] = 14'b0000101_1110100;
		logarithm_table[7697] = 14'b0000101_1110100;
		logarithm_table[7698] = 14'b0000101_1110101;
		logarithm_table[7699] = 14'b0000101_1110101;
		logarithm_table[7700] = 14'b0000101_1110101;
		logarithm_table[7701] = 14'b0000101_1110101;
		logarithm_table[7702] = 14'b0000101_1110101;
		logarithm_table[7703] = 14'b0000101_1110101;
		logarithm_table[7704] = 14'b0000101_1110101;
		logarithm_table[7705] = 14'b0000101_1110101;
		logarithm_table[7706] = 14'b0000101_1110101;
		logarithm_table[7707] = 14'b0000101_1110101;
		logarithm_table[7708] = 14'b0000101_1110101;
		logarithm_table[7709] = 14'b0000101_1110101;
		logarithm_table[7710] = 14'b0000101_1110101;
		logarithm_table[7711] = 14'b0000101_1110101;
		logarithm_table[7712] = 14'b0000101_1110101;
		logarithm_table[7713] = 14'b0000101_1110101;
		logarithm_table[7714] = 14'b0000101_1110101;
		logarithm_table[7715] = 14'b0000101_1110101;
		logarithm_table[7716] = 14'b0000101_1110101;
		logarithm_table[7717] = 14'b0000101_1110101;
		logarithm_table[7718] = 14'b0000101_1110101;
		logarithm_table[7719] = 14'b0000101_1110101;
		logarithm_table[7720] = 14'b0000101_1110101;
		logarithm_table[7721] = 14'b0000101_1110101;
		logarithm_table[7722] = 14'b0000101_1110101;
		logarithm_table[7723] = 14'b0000101_1110101;
		logarithm_table[7724] = 14'b0000101_1110101;
		logarithm_table[7725] = 14'b0000101_1110101;
		logarithm_table[7726] = 14'b0000101_1110101;
		logarithm_table[7727] = 14'b0000101_1110101;
		logarithm_table[7728] = 14'b0000101_1110101;
		logarithm_table[7729] = 14'b0000101_1110101;
		logarithm_table[7730] = 14'b0000101_1110101;
		logarithm_table[7731] = 14'b0000101_1110101;
		logarithm_table[7732] = 14'b0000101_1110101;
		logarithm_table[7733] = 14'b0000101_1110101;
		logarithm_table[7734] = 14'b0000101_1110101;
		logarithm_table[7735] = 14'b0000101_1110101;
		logarithm_table[7736] = 14'b0000101_1110101;
		logarithm_table[7737] = 14'b0000101_1110101;
		logarithm_table[7738] = 14'b0000101_1110101;
		logarithm_table[7739] = 14'b0000101_1110101;
		logarithm_table[7740] = 14'b0000101_1110110;
		logarithm_table[7741] = 14'b0000101_1110110;
		logarithm_table[7742] = 14'b0000101_1110110;
		logarithm_table[7743] = 14'b0000101_1110110;
		logarithm_table[7744] = 14'b0000101_1110110;
		logarithm_table[7745] = 14'b0000101_1110110;
		logarithm_table[7746] = 14'b0000101_1110110;
		logarithm_table[7747] = 14'b0000101_1110110;
		logarithm_table[7748] = 14'b0000101_1110110;
		logarithm_table[7749] = 14'b0000101_1110110;
		logarithm_table[7750] = 14'b0000101_1110110;
		logarithm_table[7751] = 14'b0000101_1110110;
		logarithm_table[7752] = 14'b0000101_1110110;
		logarithm_table[7753] = 14'b0000101_1110110;
		logarithm_table[7754] = 14'b0000101_1110110;
		logarithm_table[7755] = 14'b0000101_1110110;
		logarithm_table[7756] = 14'b0000101_1110110;
		logarithm_table[7757] = 14'b0000101_1110110;
		logarithm_table[7758] = 14'b0000101_1110110;
		logarithm_table[7759] = 14'b0000101_1110110;
		logarithm_table[7760] = 14'b0000101_1110110;
		logarithm_table[7761] = 14'b0000101_1110110;
		logarithm_table[7762] = 14'b0000101_1110110;
		logarithm_table[7763] = 14'b0000101_1110110;
		logarithm_table[7764] = 14'b0000101_1110110;
		logarithm_table[7765] = 14'b0000101_1110110;
		logarithm_table[7766] = 14'b0000101_1110110;
		logarithm_table[7767] = 14'b0000101_1110110;
		logarithm_table[7768] = 14'b0000101_1110110;
		logarithm_table[7769] = 14'b0000101_1110110;
		logarithm_table[7770] = 14'b0000101_1110110;
		logarithm_table[7771] = 14'b0000101_1110110;
		logarithm_table[7772] = 14'b0000101_1110110;
		logarithm_table[7773] = 14'b0000101_1110110;
		logarithm_table[7774] = 14'b0000101_1110110;
		logarithm_table[7775] = 14'b0000101_1110110;
		logarithm_table[7776] = 14'b0000101_1110110;
		logarithm_table[7777] = 14'b0000101_1110110;
		logarithm_table[7778] = 14'b0000101_1110110;
		logarithm_table[7779] = 14'b0000101_1110110;
		logarithm_table[7780] = 14'b0000101_1110110;
		logarithm_table[7781] = 14'b0000101_1110110;
		logarithm_table[7782] = 14'b0000101_1110111;
		logarithm_table[7783] = 14'b0000101_1110111;
		logarithm_table[7784] = 14'b0000101_1110111;
		logarithm_table[7785] = 14'b0000101_1110111;
		logarithm_table[7786] = 14'b0000101_1110111;
		logarithm_table[7787] = 14'b0000101_1110111;
		logarithm_table[7788] = 14'b0000101_1110111;
		logarithm_table[7789] = 14'b0000101_1110111;
		logarithm_table[7790] = 14'b0000101_1110111;
		logarithm_table[7791] = 14'b0000101_1110111;
		logarithm_table[7792] = 14'b0000101_1110111;
		logarithm_table[7793] = 14'b0000101_1110111;
		logarithm_table[7794] = 14'b0000101_1110111;
		logarithm_table[7795] = 14'b0000101_1110111;
		logarithm_table[7796] = 14'b0000101_1110111;
		logarithm_table[7797] = 14'b0000101_1110111;
		logarithm_table[7798] = 14'b0000101_1110111;
		logarithm_table[7799] = 14'b0000101_1110111;
		logarithm_table[7800] = 14'b0000101_1110111;
		logarithm_table[7801] = 14'b0000101_1110111;
		logarithm_table[7802] = 14'b0000101_1110111;
		logarithm_table[7803] = 14'b0000101_1110111;
		logarithm_table[7804] = 14'b0000101_1110111;
		logarithm_table[7805] = 14'b0000101_1110111;
		logarithm_table[7806] = 14'b0000101_1110111;
		logarithm_table[7807] = 14'b0000101_1110111;
		logarithm_table[7808] = 14'b0000101_1110111;
		logarithm_table[7809] = 14'b0000101_1110111;
		logarithm_table[7810] = 14'b0000101_1110111;
		logarithm_table[7811] = 14'b0000101_1110111;
		logarithm_table[7812] = 14'b0000101_1110111;
		logarithm_table[7813] = 14'b0000101_1110111;
		logarithm_table[7814] = 14'b0000101_1110111;
		logarithm_table[7815] = 14'b0000101_1110111;
		logarithm_table[7816] = 14'b0000101_1110111;
		logarithm_table[7817] = 14'b0000101_1110111;
		logarithm_table[7818] = 14'b0000101_1110111;
		logarithm_table[7819] = 14'b0000101_1110111;
		logarithm_table[7820] = 14'b0000101_1110111;
		logarithm_table[7821] = 14'b0000101_1110111;
		logarithm_table[7822] = 14'b0000101_1110111;
		logarithm_table[7823] = 14'b0000101_1110111;
		logarithm_table[7824] = 14'b0000101_1111000;
		logarithm_table[7825] = 14'b0000101_1111000;
		logarithm_table[7826] = 14'b0000101_1111000;
		logarithm_table[7827] = 14'b0000101_1111000;
		logarithm_table[7828] = 14'b0000101_1111000;
		logarithm_table[7829] = 14'b0000101_1111000;
		logarithm_table[7830] = 14'b0000101_1111000;
		logarithm_table[7831] = 14'b0000101_1111000;
		logarithm_table[7832] = 14'b0000101_1111000;
		logarithm_table[7833] = 14'b0000101_1111000;
		logarithm_table[7834] = 14'b0000101_1111000;
		logarithm_table[7835] = 14'b0000101_1111000;
		logarithm_table[7836] = 14'b0000101_1111000;
		logarithm_table[7837] = 14'b0000101_1111000;
		logarithm_table[7838] = 14'b0000101_1111000;
		logarithm_table[7839] = 14'b0000101_1111000;
		logarithm_table[7840] = 14'b0000101_1111000;
		logarithm_table[7841] = 14'b0000101_1111000;
		logarithm_table[7842] = 14'b0000101_1111000;
		logarithm_table[7843] = 14'b0000101_1111000;
		logarithm_table[7844] = 14'b0000101_1111000;
		logarithm_table[7845] = 14'b0000101_1111000;
		logarithm_table[7846] = 14'b0000101_1111000;
		logarithm_table[7847] = 14'b0000101_1111000;
		logarithm_table[7848] = 14'b0000101_1111000;
		logarithm_table[7849] = 14'b0000101_1111000;
		logarithm_table[7850] = 14'b0000101_1111000;
		logarithm_table[7851] = 14'b0000101_1111000;
		logarithm_table[7852] = 14'b0000101_1111000;
		logarithm_table[7853] = 14'b0000101_1111000;
		logarithm_table[7854] = 14'b0000101_1111000;
		logarithm_table[7855] = 14'b0000101_1111000;
		logarithm_table[7856] = 14'b0000101_1111000;
		logarithm_table[7857] = 14'b0000101_1111000;
		logarithm_table[7858] = 14'b0000101_1111000;
		logarithm_table[7859] = 14'b0000101_1111000;
		logarithm_table[7860] = 14'b0000101_1111000;
		logarithm_table[7861] = 14'b0000101_1111000;
		logarithm_table[7862] = 14'b0000101_1111000;
		logarithm_table[7863] = 14'b0000101_1111000;
		logarithm_table[7864] = 14'b0000101_1111000;
		logarithm_table[7865] = 14'b0000101_1111000;
		logarithm_table[7866] = 14'b0000101_1111001;
		logarithm_table[7867] = 14'b0000101_1111001;
		logarithm_table[7868] = 14'b0000101_1111001;
		logarithm_table[7869] = 14'b0000101_1111001;
		logarithm_table[7870] = 14'b0000101_1111001;
		logarithm_table[7871] = 14'b0000101_1111001;
		logarithm_table[7872] = 14'b0000101_1111001;
		logarithm_table[7873] = 14'b0000101_1111001;
		logarithm_table[7874] = 14'b0000101_1111001;
		logarithm_table[7875] = 14'b0000101_1111001;
		logarithm_table[7876] = 14'b0000101_1111001;
		logarithm_table[7877] = 14'b0000101_1111001;
		logarithm_table[7878] = 14'b0000101_1111001;
		logarithm_table[7879] = 14'b0000101_1111001;
		logarithm_table[7880] = 14'b0000101_1111001;
		logarithm_table[7881] = 14'b0000101_1111001;
		logarithm_table[7882] = 14'b0000101_1111001;
		logarithm_table[7883] = 14'b0000101_1111001;
		logarithm_table[7884] = 14'b0000101_1111001;
		logarithm_table[7885] = 14'b0000101_1111001;
		logarithm_table[7886] = 14'b0000101_1111001;
		logarithm_table[7887] = 14'b0000101_1111001;
		logarithm_table[7888] = 14'b0000101_1111001;
		logarithm_table[7889] = 14'b0000101_1111001;
		logarithm_table[7890] = 14'b0000101_1111001;
		logarithm_table[7891] = 14'b0000101_1111001;
		logarithm_table[7892] = 14'b0000101_1111001;
		logarithm_table[7893] = 14'b0000101_1111001;
		logarithm_table[7894] = 14'b0000101_1111001;
		logarithm_table[7895] = 14'b0000101_1111001;
		logarithm_table[7896] = 14'b0000101_1111001;
		logarithm_table[7897] = 14'b0000101_1111001;
		logarithm_table[7898] = 14'b0000101_1111001;
		logarithm_table[7899] = 14'b0000101_1111001;
		logarithm_table[7900] = 14'b0000101_1111001;
		logarithm_table[7901] = 14'b0000101_1111001;
		logarithm_table[7902] = 14'b0000101_1111001;
		logarithm_table[7903] = 14'b0000101_1111001;
		logarithm_table[7904] = 14'b0000101_1111001;
		logarithm_table[7905] = 14'b0000101_1111001;
		logarithm_table[7906] = 14'b0000101_1111001;
		logarithm_table[7907] = 14'b0000101_1111001;
		logarithm_table[7908] = 14'b0000101_1111001;
		logarithm_table[7909] = 14'b0000101_1111010;
		logarithm_table[7910] = 14'b0000101_1111010;
		logarithm_table[7911] = 14'b0000101_1111010;
		logarithm_table[7912] = 14'b0000101_1111010;
		logarithm_table[7913] = 14'b0000101_1111010;
		logarithm_table[7914] = 14'b0000101_1111010;
		logarithm_table[7915] = 14'b0000101_1111010;
		logarithm_table[7916] = 14'b0000101_1111010;
		logarithm_table[7917] = 14'b0000101_1111010;
		logarithm_table[7918] = 14'b0000101_1111010;
		logarithm_table[7919] = 14'b0000101_1111010;
		logarithm_table[7920] = 14'b0000101_1111010;
		logarithm_table[7921] = 14'b0000101_1111010;
		logarithm_table[7922] = 14'b0000101_1111010;
		logarithm_table[7923] = 14'b0000101_1111010;
		logarithm_table[7924] = 14'b0000101_1111010;
		logarithm_table[7925] = 14'b0000101_1111010;
		logarithm_table[7926] = 14'b0000101_1111010;
		logarithm_table[7927] = 14'b0000101_1111010;
		logarithm_table[7928] = 14'b0000101_1111010;
		logarithm_table[7929] = 14'b0000101_1111010;
		logarithm_table[7930] = 14'b0000101_1111010;
		logarithm_table[7931] = 14'b0000101_1111010;
		logarithm_table[7932] = 14'b0000101_1111010;
		logarithm_table[7933] = 14'b0000101_1111010;
		logarithm_table[7934] = 14'b0000101_1111010;
		logarithm_table[7935] = 14'b0000101_1111010;
		logarithm_table[7936] = 14'b0000101_1111010;
		logarithm_table[7937] = 14'b0000101_1111010;
		logarithm_table[7938] = 14'b0000101_1111010;
		logarithm_table[7939] = 14'b0000101_1111010;
		logarithm_table[7940] = 14'b0000101_1111010;
		logarithm_table[7941] = 14'b0000101_1111010;
		logarithm_table[7942] = 14'b0000101_1111010;
		logarithm_table[7943] = 14'b0000101_1111010;
		logarithm_table[7944] = 14'b0000101_1111010;
		logarithm_table[7945] = 14'b0000101_1111010;
		logarithm_table[7946] = 14'b0000101_1111010;
		logarithm_table[7947] = 14'b0000101_1111010;
		logarithm_table[7948] = 14'b0000101_1111010;
		logarithm_table[7949] = 14'b0000101_1111010;
		logarithm_table[7950] = 14'b0000101_1111010;
		logarithm_table[7951] = 14'b0000101_1111010;
		logarithm_table[7952] = 14'b0000101_1111011;
		logarithm_table[7953] = 14'b0000101_1111011;
		logarithm_table[7954] = 14'b0000101_1111011;
		logarithm_table[7955] = 14'b0000101_1111011;
		logarithm_table[7956] = 14'b0000101_1111011;
		logarithm_table[7957] = 14'b0000101_1111011;
		logarithm_table[7958] = 14'b0000101_1111011;
		logarithm_table[7959] = 14'b0000101_1111011;
		logarithm_table[7960] = 14'b0000101_1111011;
		logarithm_table[7961] = 14'b0000101_1111011;
		logarithm_table[7962] = 14'b0000101_1111011;
		logarithm_table[7963] = 14'b0000101_1111011;
		logarithm_table[7964] = 14'b0000101_1111011;
		logarithm_table[7965] = 14'b0000101_1111011;
		logarithm_table[7966] = 14'b0000101_1111011;
		logarithm_table[7967] = 14'b0000101_1111011;
		logarithm_table[7968] = 14'b0000101_1111011;
		logarithm_table[7969] = 14'b0000101_1111011;
		logarithm_table[7970] = 14'b0000101_1111011;
		logarithm_table[7971] = 14'b0000101_1111011;
		logarithm_table[7972] = 14'b0000101_1111011;
		logarithm_table[7973] = 14'b0000101_1111011;
		logarithm_table[7974] = 14'b0000101_1111011;
		logarithm_table[7975] = 14'b0000101_1111011;
		logarithm_table[7976] = 14'b0000101_1111011;
		logarithm_table[7977] = 14'b0000101_1111011;
		logarithm_table[7978] = 14'b0000101_1111011;
		logarithm_table[7979] = 14'b0000101_1111011;
		logarithm_table[7980] = 14'b0000101_1111011;
		logarithm_table[7981] = 14'b0000101_1111011;
		logarithm_table[7982] = 14'b0000101_1111011;
		logarithm_table[7983] = 14'b0000101_1111011;
		logarithm_table[7984] = 14'b0000101_1111011;
		logarithm_table[7985] = 14'b0000101_1111011;
		logarithm_table[7986] = 14'b0000101_1111011;
		logarithm_table[7987] = 14'b0000101_1111011;
		logarithm_table[7988] = 14'b0000101_1111011;
		logarithm_table[7989] = 14'b0000101_1111011;
		logarithm_table[7990] = 14'b0000101_1111011;
		logarithm_table[7991] = 14'b0000101_1111011;
		logarithm_table[7992] = 14'b0000101_1111011;
		logarithm_table[7993] = 14'b0000101_1111011;
		logarithm_table[7994] = 14'b0000101_1111011;
		logarithm_table[7995] = 14'b0000101_1111100;
		logarithm_table[7996] = 14'b0000101_1111100;
		logarithm_table[7997] = 14'b0000101_1111100;
		logarithm_table[7998] = 14'b0000101_1111100;
		logarithm_table[7999] = 14'b0000101_1111100;
		logarithm_table[8000] = 14'b0000101_1111100;
		logarithm_table[8001] = 14'b0000101_1111100;
		logarithm_table[8002] = 14'b0000101_1111100;
		logarithm_table[8003] = 14'b0000101_1111100;
		logarithm_table[8004] = 14'b0000101_1111100;
		logarithm_table[8005] = 14'b0000101_1111100;
		logarithm_table[8006] = 14'b0000101_1111100;
		logarithm_table[8007] = 14'b0000101_1111100;
		logarithm_table[8008] = 14'b0000101_1111100;
		logarithm_table[8009] = 14'b0000101_1111100;
		logarithm_table[8010] = 14'b0000101_1111100;
		logarithm_table[8011] = 14'b0000101_1111100;
		logarithm_table[8012] = 14'b0000101_1111100;
		logarithm_table[8013] = 14'b0000101_1111100;
		logarithm_table[8014] = 14'b0000101_1111100;
		logarithm_table[8015] = 14'b0000101_1111100;
		logarithm_table[8016] = 14'b0000101_1111100;
		logarithm_table[8017] = 14'b0000101_1111100;
		logarithm_table[8018] = 14'b0000101_1111100;
		logarithm_table[8019] = 14'b0000101_1111100;
		logarithm_table[8020] = 14'b0000101_1111100;
		logarithm_table[8021] = 14'b0000101_1111100;
		logarithm_table[8022] = 14'b0000101_1111100;
		logarithm_table[8023] = 14'b0000101_1111100;
		logarithm_table[8024] = 14'b0000101_1111100;
		logarithm_table[8025] = 14'b0000101_1111100;
		logarithm_table[8026] = 14'b0000101_1111100;
		logarithm_table[8027] = 14'b0000101_1111100;
		logarithm_table[8028] = 14'b0000101_1111100;
		logarithm_table[8029] = 14'b0000101_1111100;
		logarithm_table[8030] = 14'b0000101_1111100;
		logarithm_table[8031] = 14'b0000101_1111100;
		logarithm_table[8032] = 14'b0000101_1111100;
		logarithm_table[8033] = 14'b0000101_1111100;
		logarithm_table[8034] = 14'b0000101_1111100;
		logarithm_table[8035] = 14'b0000101_1111100;
		logarithm_table[8036] = 14'b0000101_1111100;
		logarithm_table[8037] = 14'b0000101_1111100;
		logarithm_table[8038] = 14'b0000101_1111100;
		logarithm_table[8039] = 14'b0000101_1111101;
		logarithm_table[8040] = 14'b0000101_1111101;
		logarithm_table[8041] = 14'b0000101_1111101;
		logarithm_table[8042] = 14'b0000101_1111101;
		logarithm_table[8043] = 14'b0000101_1111101;
		logarithm_table[8044] = 14'b0000101_1111101;
		logarithm_table[8045] = 14'b0000101_1111101;
		logarithm_table[8046] = 14'b0000101_1111101;
		logarithm_table[8047] = 14'b0000101_1111101;
		logarithm_table[8048] = 14'b0000101_1111101;
		logarithm_table[8049] = 14'b0000101_1111101;
		logarithm_table[8050] = 14'b0000101_1111101;
		logarithm_table[8051] = 14'b0000101_1111101;
		logarithm_table[8052] = 14'b0000101_1111101;
		logarithm_table[8053] = 14'b0000101_1111101;
		logarithm_table[8054] = 14'b0000101_1111101;
		logarithm_table[8055] = 14'b0000101_1111101;
		logarithm_table[8056] = 14'b0000101_1111101;
		logarithm_table[8057] = 14'b0000101_1111101;
		logarithm_table[8058] = 14'b0000101_1111101;
		logarithm_table[8059] = 14'b0000101_1111101;
		logarithm_table[8060] = 14'b0000101_1111101;
		logarithm_table[8061] = 14'b0000101_1111101;
		logarithm_table[8062] = 14'b0000101_1111101;
		logarithm_table[8063] = 14'b0000101_1111101;
		logarithm_table[8064] = 14'b0000101_1111101;
		logarithm_table[8065] = 14'b0000101_1111101;
		logarithm_table[8066] = 14'b0000101_1111101;
		logarithm_table[8067] = 14'b0000101_1111101;
		logarithm_table[8068] = 14'b0000101_1111101;
		logarithm_table[8069] = 14'b0000101_1111101;
		logarithm_table[8070] = 14'b0000101_1111101;
		logarithm_table[8071] = 14'b0000101_1111101;
		logarithm_table[8072] = 14'b0000101_1111101;
		logarithm_table[8073] = 14'b0000101_1111101;
		logarithm_table[8074] = 14'b0000101_1111101;
		logarithm_table[8075] = 14'b0000101_1111101;
		logarithm_table[8076] = 14'b0000101_1111101;
		logarithm_table[8077] = 14'b0000101_1111101;
		logarithm_table[8078] = 14'b0000101_1111101;
		logarithm_table[8079] = 14'b0000101_1111101;
		logarithm_table[8080] = 14'b0000101_1111101;
		logarithm_table[8081] = 14'b0000101_1111101;
		logarithm_table[8082] = 14'b0000101_1111110;
		logarithm_table[8083] = 14'b0000101_1111110;
		logarithm_table[8084] = 14'b0000101_1111110;
		logarithm_table[8085] = 14'b0000101_1111110;
		logarithm_table[8086] = 14'b0000101_1111110;
		logarithm_table[8087] = 14'b0000101_1111110;
		logarithm_table[8088] = 14'b0000101_1111110;
		logarithm_table[8089] = 14'b0000101_1111110;
		logarithm_table[8090] = 14'b0000101_1111110;
		logarithm_table[8091] = 14'b0000101_1111110;
		logarithm_table[8092] = 14'b0000101_1111110;
		logarithm_table[8093] = 14'b0000101_1111110;
		logarithm_table[8094] = 14'b0000101_1111110;
		logarithm_table[8095] = 14'b0000101_1111110;
		logarithm_table[8096] = 14'b0000101_1111110;
		logarithm_table[8097] = 14'b0000101_1111110;
		logarithm_table[8098] = 14'b0000101_1111110;
		logarithm_table[8099] = 14'b0000101_1111110;
		logarithm_table[8100] = 14'b0000101_1111110;
		logarithm_table[8101] = 14'b0000101_1111110;
		logarithm_table[8102] = 14'b0000101_1111110;
		logarithm_table[8103] = 14'b0000101_1111110;
		logarithm_table[8104] = 14'b0000101_1111110;
		logarithm_table[8105] = 14'b0000101_1111110;
		logarithm_table[8106] = 14'b0000101_1111110;
		logarithm_table[8107] = 14'b0000101_1111110;
		logarithm_table[8108] = 14'b0000101_1111110;
		logarithm_table[8109] = 14'b0000101_1111110;
		logarithm_table[8110] = 14'b0000101_1111110;
		logarithm_table[8111] = 14'b0000101_1111110;
		logarithm_table[8112] = 14'b0000101_1111110;
		logarithm_table[8113] = 14'b0000101_1111110;
		logarithm_table[8114] = 14'b0000101_1111110;
		logarithm_table[8115] = 14'b0000101_1111110;
		logarithm_table[8116] = 14'b0000101_1111110;
		logarithm_table[8117] = 14'b0000101_1111110;
		logarithm_table[8118] = 14'b0000101_1111110;
		logarithm_table[8119] = 14'b0000101_1111110;
		logarithm_table[8120] = 14'b0000101_1111110;
		logarithm_table[8121] = 14'b0000101_1111110;
		logarithm_table[8122] = 14'b0000101_1111110;
		logarithm_table[8123] = 14'b0000101_1111110;
		logarithm_table[8124] = 14'b0000101_1111110;
		logarithm_table[8125] = 14'b0000101_1111110;
		logarithm_table[8126] = 14'b0000101_1111111;
		logarithm_table[8127] = 14'b0000101_1111111;
		logarithm_table[8128] = 14'b0000101_1111111;
		logarithm_table[8129] = 14'b0000101_1111111;
		logarithm_table[8130] = 14'b0000101_1111111;
		logarithm_table[8131] = 14'b0000101_1111111;
		logarithm_table[8132] = 14'b0000101_1111111;
		logarithm_table[8133] = 14'b0000101_1111111;
		logarithm_table[8134] = 14'b0000101_1111111;
		logarithm_table[8135] = 14'b0000101_1111111;
		logarithm_table[8136] = 14'b0000101_1111111;
		logarithm_table[8137] = 14'b0000101_1111111;
		logarithm_table[8138] = 14'b0000101_1111111;
		logarithm_table[8139] = 14'b0000101_1111111;
		logarithm_table[8140] = 14'b0000101_1111111;
		logarithm_table[8141] = 14'b0000101_1111111;
		logarithm_table[8142] = 14'b0000101_1111111;
		logarithm_table[8143] = 14'b0000101_1111111;
		logarithm_table[8144] = 14'b0000101_1111111;
		logarithm_table[8145] = 14'b0000101_1111111;
		logarithm_table[8146] = 14'b0000101_1111111;
		logarithm_table[8147] = 14'b0000101_1111111;
		logarithm_table[8148] = 14'b0000101_1111111;
		logarithm_table[8149] = 14'b0000101_1111111;
		logarithm_table[8150] = 14'b0000101_1111111;
		logarithm_table[8151] = 14'b0000101_1111111;
		logarithm_table[8152] = 14'b0000101_1111111;
		logarithm_table[8153] = 14'b0000101_1111111;
		logarithm_table[8154] = 14'b0000101_1111111;
		logarithm_table[8155] = 14'b0000101_1111111;
		logarithm_table[8156] = 14'b0000101_1111111;
		logarithm_table[8157] = 14'b0000101_1111111;
		logarithm_table[8158] = 14'b0000101_1111111;
		logarithm_table[8159] = 14'b0000101_1111111;
		logarithm_table[8160] = 14'b0000101_1111111;
		logarithm_table[8161] = 14'b0000101_1111111;
		logarithm_table[8162] = 14'b0000101_1111111;
		logarithm_table[8163] = 14'b0000101_1111111;
		logarithm_table[8164] = 14'b0000101_1111111;
		logarithm_table[8165] = 14'b0000101_1111111;
		logarithm_table[8166] = 14'b0000101_1111111;
		logarithm_table[8167] = 14'b0000101_1111111;
		logarithm_table[8168] = 14'b0000101_1111111;
		logarithm_table[8169] = 14'b0000101_1111111;
		logarithm_table[8170] = 14'b0000110_0000000;
		logarithm_table[8171] = 14'b0000110_0000000;
		logarithm_table[8172] = 14'b0000110_0000000;
		logarithm_table[8173] = 14'b0000110_0000000;
		logarithm_table[8174] = 14'b0000110_0000000;
		logarithm_table[8175] = 14'b0000110_0000000;
		logarithm_table[8176] = 14'b0000110_0000000;
		logarithm_table[8177] = 14'b0000110_0000000;
		logarithm_table[8178] = 14'b0000110_0000000;
		logarithm_table[8179] = 14'b0000110_0000000;
		logarithm_table[8180] = 14'b0000110_0000000;
		logarithm_table[8181] = 14'b0000110_0000000;
		logarithm_table[8182] = 14'b0000110_0000000;
		logarithm_table[8183] = 14'b0000110_0000000;
		logarithm_table[8184] = 14'b0000110_0000000;
		logarithm_table[8185] = 14'b0000110_0000000;
		logarithm_table[8186] = 14'b0000110_0000000;
		logarithm_table[8187] = 14'b0000110_0000000;
		logarithm_table[8188] = 14'b0000110_0000000;
		logarithm_table[8189] = 14'b0000110_0000000;
		logarithm_table[8190] = 14'b0000110_0000000;
		logarithm_table[8191] = 14'b0000110_0000000;
		Dminus[1] = 14'b1111000_0111100;
		Dminus[2] = 14'b1111001_0111011;
		Dminus[3] = 14'b1111010_0000110;
		Dminus[4] = 14'b1111010_0111010;
		Dminus[5] = 14'b1111010_1100011;
		Dminus[6] = 14'b1111011_0000100;
		Dminus[7] = 14'b1111011_0100000;
		Dminus[8] = 14'b1111011_0111000;
		Dminus[9] = 14'b1111011_1001110;
		Dminus[10] = 14'b1111011_1100001;
		Dminus[11] = 14'b1111011_1110010;
		Dminus[12] = 14'b1111100_0000001;
		Dminus[13] = 14'b1111100_0010000;
		Dminus[14] = 14'b1111100_0011101;
		Dminus[15] = 14'b1111100_0101001;
		Dminus[16] = 14'b1111100_0110100;
		Dminus[17] = 14'b1111100_0111111;
		Dminus[18] = 14'b1111100_1001001;
		Dminus[19] = 14'b1111100_1010011;
		Dminus[20] = 14'b1111100_1011100;
		Dminus[21] = 14'b1111100_1100100;
		Dminus[22] = 14'b1111100_1101100;
		Dminus[23] = 14'b1111100_1110100;
		Dminus[24] = 14'b1111100_1111011;
		Dminus[25] = 14'b1111101_0000010;
		Dminus[26] = 14'b1111101_0001001;
		Dminus[27] = 14'b1111101_0010000;
		Dminus[28] = 14'b1111101_0010110;
		Dminus[29] = 14'b1111101_0011100;
		Dminus[30] = 14'b1111101_0100010;
		Dminus[31] = 14'b1111101_0100111;
		Dminus[32] = 14'b1111101_0101101;
		Dminus[33] = 14'b1111101_0110010;
		Dminus[34] = 14'b1111101_0110111;
		Dminus[35] = 14'b1111101_0111100;
		Dminus[36] = 14'b1111101_1000000;
		Dminus[37] = 14'b1111101_1000101;
		Dminus[38] = 14'b1111101_1001001;
		Dminus[39] = 14'b1111101_1001110;
		Dminus[40] = 14'b1111101_1010010;
		Dminus[41] = 14'b1111101_1010110;
		Dminus[42] = 14'b1111101_1011010;
		Dminus[43] = 14'b1111101_1011110;
		Dminus[44] = 14'b1111101_1100010;
		Dminus[45] = 14'b1111101_1100101;
		Dminus[46] = 14'b1111101_1101001;
		Dminus[47] = 14'b1111101_1101100;
		Dminus[48] = 14'b1111101_1110000;
		Dminus[49] = 14'b1111101_1110011;
		Dminus[50] = 14'b1111101_1110110;
		Dminus[51] = 14'b1111101_1111001;
		Dminus[52] = 14'b1111101_1111101;
		Dminus[53] = 14'b1111110_0000000;
		Dminus[54] = 14'b1111110_0000011;
		Dminus[55] = 14'b1111110_0000110;
		Dminus[56] = 14'b1111110_0001000;
		Dminus[57] = 14'b1111110_0001011;
		Dminus[58] = 14'b1111110_0001110;
		Dminus[59] = 14'b1111110_0010001;
		Dminus[60] = 14'b1111110_0010011;
		Dminus[61] = 14'b1111110_0010110;
		Dminus[62] = 14'b1111110_0011000;
		Dminus[63] = 14'b1111110_0011011;
		Dminus[64] = 14'b1111110_0011101;
		Dminus[65] = 14'b1111110_0100000;
		Dminus[66] = 14'b1111110_0100010;
		Dminus[67] = 14'b1111110_0100100;
		Dminus[68] = 14'b1111110_0100111;
		Dminus[69] = 14'b1111110_0101001;
		Dminus[70] = 14'b1111110_0101011;
		Dminus[71] = 14'b1111110_0101101;
		Dminus[72] = 14'b1111110_0101111;
		Dminus[73] = 14'b1111110_0110001;
		Dminus[74] = 14'b1111110_0110011;
		Dminus[75] = 14'b1111110_0110101;
		Dminus[76] = 14'b1111110_0110111;
		Dminus[77] = 14'b1111110_0111001;
		Dminus[78] = 14'b1111110_0111011;
		Dminus[79] = 14'b1111110_0111101;
		Dminus[80] = 14'b1111110_0111111;
		Dminus[81] = 14'b1111110_1000001;
		Dminus[82] = 14'b1111110_1000011;
		Dminus[83] = 14'b1111110_1000100;
		Dminus[84] = 14'b1111110_1000110;
		Dminus[85] = 14'b1111110_1001000;
		Dminus[86] = 14'b1111110_1001010;
		Dminus[87] = 14'b1111110_1001011;
		Dminus[88] = 14'b1111110_1001101;
		Dminus[89] = 14'b1111110_1001110;
		Dminus[90] = 14'b1111110_1010000;
		Dminus[91] = 14'b1111110_1010010;
		Dminus[92] = 14'b1111110_1010011;
		Dminus[93] = 14'b1111110_1010101;
		Dminus[94] = 14'b1111110_1010110;
		Dminus[95] = 14'b1111110_1011000;
		Dminus[96] = 14'b1111110_1011001;
		Dminus[97] = 14'b1111110_1011011;
		Dminus[98] = 14'b1111110_1011100;
		Dminus[99] = 14'b1111110_1011110;
		Dminus[100] = 14'b1111110_1011111;
		Dminus[101] = 14'b1111110_1100000;
		Dminus[102] = 14'b1111110_1100010;
		Dminus[103] = 14'b1111110_1100011;
		Dminus[104] = 14'b1111110_1100100;
		Dminus[105] = 14'b1111110_1100110;
		Dminus[106] = 14'b1111110_1100111;
		Dminus[107] = 14'b1111110_1101000;
		Dminus[108] = 14'b1111110_1101010;
		Dminus[109] = 14'b1111110_1101011;
		Dminus[110] = 14'b1111110_1101100;
		Dminus[111] = 14'b1111110_1101101;
		Dminus[112] = 14'b1111110_1101110;
		Dminus[113] = 14'b1111110_1110000;
		Dminus[114] = 14'b1111110_1110001;
		Dminus[115] = 14'b1111110_1110010;
		Dminus[116] = 14'b1111110_1110011;
		Dminus[117] = 14'b1111110_1110100;
		Dminus[118] = 14'b1111110_1110101;
		Dminus[119] = 14'b1111110_1110111;
		Dminus[120] = 14'b1111110_1111000;
		Dminus[121] = 14'b1111110_1111001;
		Dminus[122] = 14'b1111110_1111010;
		Dminus[123] = 14'b1111110_1111011;
		Dminus[124] = 14'b1111110_1111100;
		Dminus[125] = 14'b1111110_1111101;
		Dminus[126] = 14'b1111110_1111110;
		Dminus[127] = 14'b1111110_1111111;
		Dminus[128] = 14'b1111111_0000000;
		Dminus[129] = 14'b1111111_0000001;
		Dminus[130] = 14'b1111111_0000010;
		Dminus[131] = 14'b1111111_0000011;
		Dminus[132] = 14'b1111111_0000100;
		Dminus[133] = 14'b1111111_0000101;
		Dminus[134] = 14'b1111111_0000110;
		Dminus[135] = 14'b1111111_0000111;
		Dminus[136] = 14'b1111111_0001000;
		Dminus[137] = 14'b1111111_0001001;
		Dminus[138] = 14'b1111111_0001001;
		Dminus[139] = 14'b1111111_0001010;
		Dminus[140] = 14'b1111111_0001011;
		Dminus[141] = 14'b1111111_0001100;
		Dminus[142] = 14'b1111111_0001101;
		Dminus[143] = 14'b1111111_0001110;
		Dminus[144] = 14'b1111111_0001111;
		Dminus[145] = 14'b1111111_0010000;
		Dminus[146] = 14'b1111111_0010000;
		Dminus[147] = 14'b1111111_0010001;
		Dminus[148] = 14'b1111111_0010010;
		Dminus[149] = 14'b1111111_0010011;
		Dminus[150] = 14'b1111111_0010100;
		Dminus[151] = 14'b1111111_0010100;
		Dminus[152] = 14'b1111111_0010101;
		Dminus[153] = 14'b1111111_0010110;
		Dminus[154] = 14'b1111111_0010111;
		Dminus[155] = 14'b1111111_0011000;
		Dminus[156] = 14'b1111111_0011000;
		Dminus[157] = 14'b1111111_0011001;
		Dminus[158] = 14'b1111111_0011010;
		Dminus[159] = 14'b1111111_0011011;
		Dminus[160] = 14'b1111111_0011011;
		Dminus[161] = 14'b1111111_0011100;
		Dminus[162] = 14'b1111111_0011101;
		Dminus[163] = 14'b1111111_0011101;
		Dminus[164] = 14'b1111111_0011110;
		Dminus[165] = 14'b1111111_0011111;
		Dminus[166] = 14'b1111111_0011111;
		Dminus[167] = 14'b1111111_0100000;
		Dminus[168] = 14'b1111111_0100001;
		Dminus[169] = 14'b1111111_0100010;
		Dminus[170] = 14'b1111111_0100010;
		Dminus[171] = 14'b1111111_0100011;
		Dminus[172] = 14'b1111111_0100100;
		Dminus[173] = 14'b1111111_0100100;
		Dminus[174] = 14'b1111111_0100101;
		Dminus[175] = 14'b1111111_0100101;
		Dminus[176] = 14'b1111111_0100110;
		Dminus[177] = 14'b1111111_0100111;
		Dminus[178] = 14'b1111111_0100111;
		Dminus[179] = 14'b1111111_0101000;
		Dminus[180] = 14'b1111111_0101001;
		Dminus[181] = 14'b1111111_0101001;
		Dminus[182] = 14'b1111111_0101010;
		Dminus[183] = 14'b1111111_0101010;
		Dminus[184] = 14'b1111111_0101011;
		Dminus[185] = 14'b1111111_0101011;
		Dminus[186] = 14'b1111111_0101100;
		Dminus[187] = 14'b1111111_0101101;
		Dminus[188] = 14'b1111111_0101101;
		Dminus[189] = 14'b1111111_0101110;
		Dminus[190] = 14'b1111111_0101110;
		Dminus[191] = 14'b1111111_0101111;
		Dminus[192] = 14'b1111111_0101111;
		Dminus[193] = 14'b1111111_0110000;
		Dminus[194] = 14'b1111111_0110001;
		Dminus[195] = 14'b1111111_0110001;
		Dminus[196] = 14'b1111111_0110010;
		Dminus[197] = 14'b1111111_0110010;
		Dminus[198] = 14'b1111111_0110011;
		Dminus[199] = 14'b1111111_0110011;
		Dminus[200] = 14'b1111111_0110100;
		Dminus[201] = 14'b1111111_0110100;
		Dminus[202] = 14'b1111111_0110101;
		Dminus[203] = 14'b1111111_0110101;
		Dminus[204] = 14'b1111111_0110110;
		Dminus[205] = 14'b1111111_0110110;
		Dminus[206] = 14'b1111111_0110111;
		Dminus[207] = 14'b1111111_0110111;
		Dminus[208] = 14'b1111111_0111000;
		Dminus[209] = 14'b1111111_0111000;
		Dminus[210] = 14'b1111111_0111001;
		Dminus[211] = 14'b1111111_0111001;
		Dminus[212] = 14'b1111111_0111010;
		Dminus[213] = 14'b1111111_0111010;
		Dminus[214] = 14'b1111111_0111010;
		Dminus[215] = 14'b1111111_0111011;
		Dminus[216] = 14'b1111111_0111011;
		Dminus[217] = 14'b1111111_0111100;
		Dminus[218] = 14'b1111111_0111100;
		Dminus[219] = 14'b1111111_0111101;
		Dminus[220] = 14'b1111111_0111101;
		Dminus[221] = 14'b1111111_0111110;
		Dminus[222] = 14'b1111111_0111110;
		Dminus[223] = 14'b1111111_0111110;
		Dminus[224] = 14'b1111111_0111111;
		Dminus[225] = 14'b1111111_0111111;
		Dminus[226] = 14'b1111111_1000000;
		Dminus[227] = 14'b1111111_1000000;
		Dminus[228] = 14'b1111111_1000001;
		Dminus[229] = 14'b1111111_1000001;
		Dminus[230] = 14'b1111111_1000001;
		Dminus[231] = 14'b1111111_1000010;
		Dminus[232] = 14'b1111111_1000010;
		Dminus[233] = 14'b1111111_1000011;
		Dminus[234] = 14'b1111111_1000011;
		Dminus[235] = 14'b1111111_1000011;
		Dminus[236] = 14'b1111111_1000100;
		Dminus[237] = 14'b1111111_1000100;
		Dminus[238] = 14'b1111111_1000100;
		Dminus[239] = 14'b1111111_1000101;
		Dminus[240] = 14'b1111111_1000101;
		Dminus[241] = 14'b1111111_1000110;
		Dminus[242] = 14'b1111111_1000110;
		Dminus[243] = 14'b1111111_1000110;
		Dminus[244] = 14'b1111111_1000111;
		Dminus[245] = 14'b1111111_1000111;
		Dminus[246] = 14'b1111111_1000111;
		Dminus[247] = 14'b1111111_1001000;
		Dminus[248] = 14'b1111111_1001000;
		Dminus[249] = 14'b1111111_1001000;
		Dminus[250] = 14'b1111111_1001001;
		Dminus[251] = 14'b1111111_1001001;
		Dminus[252] = 14'b1111111_1001010;
		Dminus[253] = 14'b1111111_1001010;
		Dminus[254] = 14'b1111111_1001010;
		Dminus[255] = 14'b1111111_1001011;
		Dminus[256] = 14'b1111111_1001011;
		Dminus[257] = 14'b1111111_1001011;
		Dminus[258] = 14'b1111111_1001100;
		Dminus[259] = 14'b1111111_1001100;
		Dminus[260] = 14'b1111111_1001100;
		Dminus[261] = 14'b1111111_1001101;
		Dminus[262] = 14'b1111111_1001101;
		Dminus[263] = 14'b1111111_1001101;
		Dminus[264] = 14'b1111111_1001101;
		Dminus[265] = 14'b1111111_1001110;
		Dminus[266] = 14'b1111111_1001110;
		Dminus[267] = 14'b1111111_1001110;
		Dminus[268] = 14'b1111111_1001111;
		Dminus[269] = 14'b1111111_1001111;
		Dminus[270] = 14'b1111111_1001111;
		Dminus[271] = 14'b1111111_1010000;
		Dminus[272] = 14'b1111111_1010000;
		Dminus[273] = 14'b1111111_1010000;
		Dminus[274] = 14'b1111111_1010001;
		Dminus[275] = 14'b1111111_1010001;
		Dminus[276] = 14'b1111111_1010001;
		Dminus[277] = 14'b1111111_1010001;
		Dminus[278] = 14'b1111111_1010010;
		Dminus[279] = 14'b1111111_1010010;
		Dminus[280] = 14'b1111111_1010010;
		Dminus[281] = 14'b1111111_1010011;
		Dminus[282] = 14'b1111111_1010011;
		Dminus[283] = 14'b1111111_1010011;
		Dminus[284] = 14'b1111111_1010011;
		Dminus[285] = 14'b1111111_1010100;
		Dminus[286] = 14'b1111111_1010100;
		Dminus[287] = 14'b1111111_1010100;
		Dminus[288] = 14'b1111111_1010100;
		Dminus[289] = 14'b1111111_1010101;
		Dminus[290] = 14'b1111111_1010101;
		Dminus[291] = 14'b1111111_1010101;
		Dminus[292] = 14'b1111111_1010101;
		Dminus[293] = 14'b1111111_1010110;
		Dminus[294] = 14'b1111111_1010110;
		Dminus[295] = 14'b1111111_1010110;
		Dminus[296] = 14'b1111111_1010110;
		Dminus[297] = 14'b1111111_1010111;
		Dminus[298] = 14'b1111111_1010111;
		Dminus[299] = 14'b1111111_1010111;
		Dminus[300] = 14'b1111111_1010111;
		Dminus[301] = 14'b1111111_1011000;
		Dminus[302] = 14'b1111111_1011000;
		Dminus[303] = 14'b1111111_1011000;
		Dminus[304] = 14'b1111111_1011000;
		Dminus[305] = 14'b1111111_1011001;
		Dminus[306] = 14'b1111111_1011001;
		Dminus[307] = 14'b1111111_1011001;
		Dminus[308] = 14'b1111111_1011001;
		Dminus[309] = 14'b1111111_1011010;
		Dminus[310] = 14'b1111111_1011010;
		Dminus[311] = 14'b1111111_1011010;
		Dminus[312] = 14'b1111111_1011010;
		Dminus[313] = 14'b1111111_1011011;
		Dminus[314] = 14'b1111111_1011011;
		Dminus[315] = 14'b1111111_1011011;
		Dminus[316] = 14'b1111111_1011011;
		Dminus[317] = 14'b1111111_1011011;
		Dminus[318] = 14'b1111111_1011100;
		Dminus[319] = 14'b1111111_1011100;
		Dminus[320] = 14'b1111111_1011100;
		Dminus[321] = 14'b1111111_1011100;
		Dminus[322] = 14'b1111111_1011101;
		Dminus[323] = 14'b1111111_1011101;
		Dminus[324] = 14'b1111111_1011101;
		Dminus[325] = 14'b1111111_1011101;
		Dminus[326] = 14'b1111111_1011101;
		Dminus[327] = 14'b1111111_1011110;
		Dminus[328] = 14'b1111111_1011110;
		Dminus[329] = 14'b1111111_1011110;
		Dminus[330] = 14'b1111111_1011110;
		Dminus[331] = 14'b1111111_1011110;
		Dminus[332] = 14'b1111111_1011111;
		Dminus[333] = 14'b1111111_1011111;
		Dminus[334] = 14'b1111111_1011111;
		Dminus[335] = 14'b1111111_1011111;
		Dminus[336] = 14'b1111111_1011111;
		Dminus[337] = 14'b1111111_1100000;
		Dminus[338] = 14'b1111111_1100000;
		Dminus[339] = 14'b1111111_1100000;
		Dminus[340] = 14'b1111111_1100000;
		Dminus[341] = 14'b1111111_1100000;
		Dminus[342] = 14'b1111111_1100000;
		Dminus[343] = 14'b1111111_1100001;
		Dminus[344] = 14'b1111111_1100001;
		Dminus[345] = 14'b1111111_1100001;
		Dminus[346] = 14'b1111111_1100001;
		Dminus[347] = 14'b1111111_1100001;
		Dminus[348] = 14'b1111111_1100010;
		Dminus[349] = 14'b1111111_1100010;
		Dminus[350] = 14'b1111111_1100010;
		Dminus[351] = 14'b1111111_1100010;
		Dminus[352] = 14'b1111111_1100010;
		Dminus[353] = 14'b1111111_1100010;
		Dminus[354] = 14'b1111111_1100011;
		Dminus[355] = 14'b1111111_1100011;
		Dminus[356] = 14'b1111111_1100011;
		Dminus[357] = 14'b1111111_1100011;
		Dminus[358] = 14'b1111111_1100011;
		Dminus[359] = 14'b1111111_1100011;
		Dminus[360] = 14'b1111111_1100100;
		Dminus[361] = 14'b1111111_1100100;
		Dminus[362] = 14'b1111111_1100100;
		Dminus[363] = 14'b1111111_1100100;
		Dminus[364] = 14'b1111111_1100100;
		Dminus[365] = 14'b1111111_1100100;
		Dminus[366] = 14'b1111111_1100101;
		Dminus[367] = 14'b1111111_1100101;
		Dminus[368] = 14'b1111111_1100101;
		Dminus[369] = 14'b1111111_1100101;
		Dminus[370] = 14'b1111111_1100101;
		Dminus[371] = 14'b1111111_1100101;
		Dminus[372] = 14'b1111111_1100110;
		Dminus[373] = 14'b1111111_1100110;
		Dminus[374] = 14'b1111111_1100110;
		Dminus[375] = 14'b1111111_1100110;
		Dminus[376] = 14'b1111111_1100110;
		Dminus[377] = 14'b1111111_1100110;
		Dminus[378] = 14'b1111111_1100110;
		Dminus[379] = 14'b1111111_1100111;
		Dminus[380] = 14'b1111111_1100111;
		Dminus[381] = 14'b1111111_1100111;
		Dminus[382] = 14'b1111111_1100111;
		Dminus[383] = 14'b1111111_1100111;
		Dminus[384] = 14'b1111111_1100111;
		Dminus[385] = 14'b1111111_1100111;
		Dminus[386] = 14'b1111111_1101000;
		Dminus[387] = 14'b1111111_1101000;
		Dminus[388] = 14'b1111111_1101000;
		Dminus[389] = 14'b1111111_1101000;
		Dminus[390] = 14'b1111111_1101000;
		Dminus[391] = 14'b1111111_1101000;
		Dminus[392] = 14'b1111111_1101000;
		Dminus[393] = 14'b1111111_1101001;
		Dminus[394] = 14'b1111111_1101001;
		Dminus[395] = 14'b1111111_1101001;
		Dminus[396] = 14'b1111111_1101001;
		Dminus[397] = 14'b1111111_1101001;
		Dminus[398] = 14'b1111111_1101001;
		Dminus[399] = 14'b1111111_1101001;
		Dminus[400] = 14'b1111111_1101010;
		Dminus[401] = 14'b1111111_1101010;
		Dminus[402] = 14'b1111111_1101010;
		Dminus[403] = 14'b1111111_1101010;
		Dminus[404] = 14'b1111111_1101010;
		Dminus[405] = 14'b1111111_1101010;
		Dminus[406] = 14'b1111111_1101010;
		Dminus[407] = 14'b1111111_1101010;
		Dminus[408] = 14'b1111111_1101011;
		Dminus[409] = 14'b1111111_1101011;
		Dminus[410] = 14'b1111111_1101011;
		Dminus[411] = 14'b1111111_1101011;
		Dminus[412] = 14'b1111111_1101011;
		Dminus[413] = 14'b1111111_1101011;
		Dminus[414] = 14'b1111111_1101011;
		Dminus[415] = 14'b1111111_1101011;
		Dminus[416] = 14'b1111111_1101011;
		Dminus[417] = 14'b1111111_1101100;
		Dminus[418] = 14'b1111111_1101100;
		Dminus[419] = 14'b1111111_1101100;
		Dminus[420] = 14'b1111111_1101100;
		Dminus[421] = 14'b1111111_1101100;
		Dminus[422] = 14'b1111111_1101100;
		Dminus[423] = 14'b1111111_1101100;
		Dminus[424] = 14'b1111111_1101100;
		Dminus[425] = 14'b1111111_1101101;
		Dminus[426] = 14'b1111111_1101101;
		Dminus[427] = 14'b1111111_1101101;
		Dminus[428] = 14'b1111111_1101101;
		Dminus[429] = 14'b1111111_1101101;
		Dminus[430] = 14'b1111111_1101101;
		Dminus[431] = 14'b1111111_1101101;
		Dminus[432] = 14'b1111111_1101101;
		Dminus[433] = 14'b1111111_1101101;
		Dminus[434] = 14'b1111111_1101101;
		Dminus[435] = 14'b1111111_1101110;
		Dminus[436] = 14'b1111111_1101110;
		Dminus[437] = 14'b1111111_1101110;
		Dminus[438] = 14'b1111111_1101110;
		Dminus[439] = 14'b1111111_1101110;
		Dminus[440] = 14'b1111111_1101110;
		Dminus[441] = 14'b1111111_1101110;
		Dminus[442] = 14'b1111111_1101110;
		Dminus[443] = 14'b1111111_1101110;
		Dminus[444] = 14'b1111111_1101111;
		Dminus[445] = 14'b1111111_1101111;
		Dminus[446] = 14'b1111111_1101111;
		Dminus[447] = 14'b1111111_1101111;
		Dminus[448] = 14'b1111111_1101111;
		Dminus[449] = 14'b1111111_1101111;
		Dminus[450] = 14'b1111111_1101111;
		Dminus[451] = 14'b1111111_1101111;
		Dminus[452] = 14'b1111111_1101111;
		Dminus[453] = 14'b1111111_1101111;
		Dminus[454] = 14'b1111111_1101111;
		Dminus[455] = 14'b1111111_1110000;
		Dminus[456] = 14'b1111111_1110000;
		Dminus[457] = 14'b1111111_1110000;
		Dminus[458] = 14'b1111111_1110000;
		Dminus[459] = 14'b1111111_1110000;
		Dminus[460] = 14'b1111111_1110000;
		Dminus[461] = 14'b1111111_1110000;
		Dminus[462] = 14'b1111111_1110000;
		Dminus[463] = 14'b1111111_1110000;
		Dminus[464] = 14'b1111111_1110000;
		Dminus[465] = 14'b1111111_1110000;
		Dminus[466] = 14'b1111111_1110001;
		Dminus[467] = 14'b1111111_1110001;
		Dminus[468] = 14'b1111111_1110001;
		Dminus[469] = 14'b1111111_1110001;
		Dminus[470] = 14'b1111111_1110001;
		Dminus[471] = 14'b1111111_1110001;
		Dminus[472] = 14'b1111111_1110001;
		Dminus[473] = 14'b1111111_1110001;
		Dminus[474] = 14'b1111111_1110001;
		Dminus[475] = 14'b1111111_1110001;
		Dminus[476] = 14'b1111111_1110001;
		Dminus[477] = 14'b1111111_1110001;
		Dminus[478] = 14'b1111111_1110010;
		Dminus[479] = 14'b1111111_1110010;
		Dminus[480] = 14'b1111111_1110010;
		Dminus[481] = 14'b1111111_1110010;
		Dminus[482] = 14'b1111111_1110010;
		Dminus[483] = 14'b1111111_1110010;
		Dminus[484] = 14'b1111111_1110010;
		Dminus[485] = 14'b1111111_1110010;
		Dminus[486] = 14'b1111111_1110010;
		Dminus[487] = 14'b1111111_1110010;
		Dminus[488] = 14'b1111111_1110010;
		Dminus[489] = 14'b1111111_1110010;
		Dminus[490] = 14'b1111111_1110011;
		Dminus[491] = 14'b1111111_1110011;
		Dminus[492] = 14'b1111111_1110011;
		Dminus[493] = 14'b1111111_1110011;
		Dminus[494] = 14'b1111111_1110011;
		Dminus[495] = 14'b1111111_1110011;
		Dminus[496] = 14'b1111111_1110011;
		Dminus[497] = 14'b1111111_1110011;
		Dminus[498] = 14'b1111111_1110011;
		Dminus[499] = 14'b1111111_1110011;
		Dminus[500] = 14'b1111111_1110011;
		Dminus[501] = 14'b1111111_1110011;
		Dminus[502] = 14'b1111111_1110011;
		Dminus[503] = 14'b1111111_1110011;
		Dminus[504] = 14'b1111111_1110100;
		Dminus[505] = 14'b1111111_1110100;
		Dminus[506] = 14'b1111111_1110100;
		Dminus[507] = 14'b1111111_1110100;
		Dminus[508] = 14'b1111111_1110100;
		Dminus[509] = 14'b1111111_1110100;
		Dminus[510] = 14'b1111111_1110100;
		Dminus[511] = 14'b1111111_1110100;
		Dminus[512] = 14'b1111111_1110100;
		Dminus[513] = 14'b1111111_1110100;
		Dminus[514] = 14'b1111111_1110100;
		Dminus[515] = 14'b1111111_1110100;
		Dminus[516] = 14'b1111111_1110100;
		Dminus[517] = 14'b1111111_1110100;
		Dminus[518] = 14'b1111111_1110100;
		Dminus[519] = 14'b1111111_1110101;
		Dminus[520] = 14'b1111111_1110101;
		Dminus[521] = 14'b1111111_1110101;
		Dminus[522] = 14'b1111111_1110101;
		Dminus[523] = 14'b1111111_1110101;
		Dminus[524] = 14'b1111111_1110101;
		Dminus[525] = 14'b1111111_1110101;
		Dminus[526] = 14'b1111111_1110101;
		Dminus[527] = 14'b1111111_1110101;
		Dminus[528] = 14'b1111111_1110101;
		Dminus[529] = 14'b1111111_1110101;
		Dminus[530] = 14'b1111111_1110101;
		Dminus[531] = 14'b1111111_1110101;
		Dminus[532] = 14'b1111111_1110101;
		Dminus[533] = 14'b1111111_1110101;
		Dminus[534] = 14'b1111111_1110101;
		Dminus[535] = 14'b1111111_1110110;
		Dminus[536] = 14'b1111111_1110110;
		Dminus[537] = 14'b1111111_1110110;
		Dminus[538] = 14'b1111111_1110110;
		Dminus[539] = 14'b1111111_1110110;
		Dminus[540] = 14'b1111111_1110110;
		Dminus[541] = 14'b1111111_1110110;
		Dminus[542] = 14'b1111111_1110110;
		Dminus[543] = 14'b1111111_1110110;
		Dminus[544] = 14'b1111111_1110110;
		Dminus[545] = 14'b1111111_1110110;
		Dminus[546] = 14'b1111111_1110110;
		Dminus[547] = 14'b1111111_1110110;
		Dminus[548] = 14'b1111111_1110110;
		Dminus[549] = 14'b1111111_1110110;
		Dminus[550] = 14'b1111111_1110110;
		Dminus[551] = 14'b1111111_1110110;
		Dminus[552] = 14'b1111111_1110110;
		Dminus[553] = 14'b1111111_1110111;
		Dminus[554] = 14'b1111111_1110111;
		Dminus[555] = 14'b1111111_1110111;
		Dminus[556] = 14'b1111111_1110111;
		Dminus[557] = 14'b1111111_1110111;
		Dminus[558] = 14'b1111111_1110111;
		Dminus[559] = 14'b1111111_1110111;
		Dminus[560] = 14'b1111111_1110111;
		Dminus[561] = 14'b1111111_1110111;
		Dminus[562] = 14'b1111111_1110111;
		Dminus[563] = 14'b1111111_1110111;
		Dminus[564] = 14'b1111111_1110111;
		Dminus[565] = 14'b1111111_1110111;
		Dminus[566] = 14'b1111111_1110111;
		Dminus[567] = 14'b1111111_1110111;
		Dminus[568] = 14'b1111111_1110111;
		Dminus[569] = 14'b1111111_1110111;
		Dminus[570] = 14'b1111111_1110111;
		Dminus[571] = 14'b1111111_1110111;
		Dminus[572] = 14'b1111111_1110111;
		Dminus[573] = 14'b1111111_1111000;
		Dminus[574] = 14'b1111111_1111000;
		Dminus[575] = 14'b1111111_1111000;
		Dminus[576] = 14'b1111111_1111000;
		Dminus[577] = 14'b1111111_1111000;
		Dminus[578] = 14'b1111111_1111000;
		Dminus[579] = 14'b1111111_1111000;
		Dminus[580] = 14'b1111111_1111000;
		Dminus[581] = 14'b1111111_1111000;
		Dminus[582] = 14'b1111111_1111000;
		Dminus[583] = 14'b1111111_1111000;
		Dminus[584] = 14'b1111111_1111000;
		Dminus[585] = 14'b1111111_1111000;
		Dminus[586] = 14'b1111111_1111000;
		Dminus[587] = 14'b1111111_1111000;
		Dminus[588] = 14'b1111111_1111000;
		Dminus[589] = 14'b1111111_1111000;
		Dminus[590] = 14'b1111111_1111000;
		Dminus[591] = 14'b1111111_1111000;
		Dminus[592] = 14'b1111111_1111000;
		Dminus[593] = 14'b1111111_1111000;
		Dminus[594] = 14'b1111111_1111000;
		Dminus[595] = 14'b1111111_1111000;
		Dminus[596] = 14'b1111111_1111001;
		Dminus[597] = 14'b1111111_1111001;
		Dminus[598] = 14'b1111111_1111001;
		Dminus[599] = 14'b1111111_1111001;
		Dminus[600] = 14'b1111111_1111001;
		Dminus[601] = 14'b1111111_1111001;
		Dminus[602] = 14'b1111111_1111001;
		Dminus[603] = 14'b1111111_1111001;
		Dminus[604] = 14'b1111111_1111001;
		Dminus[605] = 14'b1111111_1111001;
		Dminus[606] = 14'b1111111_1111001;
		Dminus[607] = 14'b1111111_1111001;
		Dminus[608] = 14'b1111111_1111001;
		Dminus[609] = 14'b1111111_1111001;
		Dminus[610] = 14'b1111111_1111001;
		Dminus[611] = 14'b1111111_1111001;
		Dminus[612] = 14'b1111111_1111001;
		Dminus[613] = 14'b1111111_1111001;
		Dminus[614] = 14'b1111111_1111001;
		Dminus[615] = 14'b1111111_1111001;
		Dminus[616] = 14'b1111111_1111001;
		Dminus[617] = 14'b1111111_1111001;
		Dminus[618] = 14'b1111111_1111001;
		Dminus[619] = 14'b1111111_1111001;
		Dminus[620] = 14'b1111111_1111001;
		Dminus[621] = 14'b1111111_1111001;
		Dminus[622] = 14'b1111111_1111010;
		Dminus[623] = 14'b1111111_1111010;
		Dminus[624] = 14'b1111111_1111010;
		Dminus[625] = 14'b1111111_1111010;
		Dminus[626] = 14'b1111111_1111010;
		Dminus[627] = 14'b1111111_1111010;
		Dminus[628] = 14'b1111111_1111010;
		Dminus[629] = 14'b1111111_1111010;
		Dminus[630] = 14'b1111111_1111010;
		Dminus[631] = 14'b1111111_1111010;
		Dminus[632] = 14'b1111111_1111010;
		Dminus[633] = 14'b1111111_1111010;
		Dminus[634] = 14'b1111111_1111010;
		Dminus[635] = 14'b1111111_1111010;
		Dminus[636] = 14'b1111111_1111010;
		Dminus[637] = 14'b1111111_1111010;
		Dminus[638] = 14'b1111111_1111010;
		Dminus[639] = 14'b1111111_1111010;
		Dminus[640] = 14'b1111111_1111010;
		Dminus[641] = 14'b1111111_1111010;
		Dminus[642] = 14'b1111111_1111010;
		Dminus[643] = 14'b1111111_1111010;
		Dminus[644] = 14'b1111111_1111010;
		Dminus[645] = 14'b1111111_1111010;
		Dminus[646] = 14'b1111111_1111010;
		Dminus[647] = 14'b1111111_1111010;
		Dminus[648] = 14'b1111111_1111010;
		Dminus[649] = 14'b1111111_1111010;
		Dminus[650] = 14'b1111111_1111010;
		Dminus[651] = 14'b1111111_1111010;
		Dminus[652] = 14'b1111111_1111011;
		Dminus[653] = 14'b1111111_1111011;
		Dminus[654] = 14'b1111111_1111011;
		Dminus[655] = 14'b1111111_1111011;
		Dminus[656] = 14'b1111111_1111011;
		Dminus[657] = 14'b1111111_1111011;
		Dminus[658] = 14'b1111111_1111011;
		Dminus[659] = 14'b1111111_1111011;
		Dminus[660] = 14'b1111111_1111011;
		Dminus[661] = 14'b1111111_1111011;
		Dminus[662] = 14'b1111111_1111011;
		Dminus[663] = 14'b1111111_1111011;
		Dminus[664] = 14'b1111111_1111011;
		Dminus[665] = 14'b1111111_1111011;
		Dminus[666] = 14'b1111111_1111011;
		Dminus[667] = 14'b1111111_1111011;
		Dminus[668] = 14'b1111111_1111011;
		Dminus[669] = 14'b1111111_1111011;
		Dminus[670] = 14'b1111111_1111011;
		Dminus[671] = 14'b1111111_1111011;
		Dminus[672] = 14'b1111111_1111011;
		Dminus[673] = 14'b1111111_1111011;
		Dminus[674] = 14'b1111111_1111011;
		Dminus[675] = 14'b1111111_1111011;
		Dminus[676] = 14'b1111111_1111011;
		Dminus[677] = 14'b1111111_1111011;
		Dminus[678] = 14'b1111111_1111011;
		Dminus[679] = 14'b1111111_1111011;
		Dminus[680] = 14'b1111111_1111011;
		Dminus[681] = 14'b1111111_1111011;
		Dminus[682] = 14'b1111111_1111011;
		Dminus[683] = 14'b1111111_1111011;
		Dminus[684] = 14'b1111111_1111011;
		Dminus[685] = 14'b1111111_1111011;
		Dminus[686] = 14'b1111111_1111011;
		Dminus[687] = 14'b1111111_1111011;
		Dminus[688] = 14'b1111111_1111011;
		Dminus[689] = 14'b1111111_1111100;
		Dminus[690] = 14'b1111111_1111100;
		Dminus[691] = 14'b1111111_1111100;
		Dminus[692] = 14'b1111111_1111100;
		Dminus[693] = 14'b1111111_1111100;
		Dminus[694] = 14'b1111111_1111100;
		Dminus[695] = 14'b1111111_1111100;
		Dminus[696] = 14'b1111111_1111100;
		Dminus[697] = 14'b1111111_1111100;
		Dminus[698] = 14'b1111111_1111100;
		Dminus[699] = 14'b1111111_1111100;
		Dminus[700] = 14'b1111111_1111100;
		Dminus[701] = 14'b1111111_1111100;
		Dminus[702] = 14'b1111111_1111100;
		Dminus[703] = 14'b1111111_1111100;
		Dminus[704] = 14'b1111111_1111100;
		Dminus[705] = 14'b1111111_1111100;
		Dminus[706] = 14'b1111111_1111100;
		Dminus[707] = 14'b1111111_1111100;
		Dminus[708] = 14'b1111111_1111100;
		Dminus[709] = 14'b1111111_1111100;
		Dminus[710] = 14'b1111111_1111100;
		Dminus[711] = 14'b1111111_1111100;
		Dminus[712] = 14'b1111111_1111100;
		Dminus[713] = 14'b1111111_1111100;
		Dminus[714] = 14'b1111111_1111100;
		Dminus[715] = 14'b1111111_1111100;
		Dminus[716] = 14'b1111111_1111100;
		Dminus[717] = 14'b1111111_1111100;
		Dminus[718] = 14'b1111111_1111100;
		Dminus[719] = 14'b1111111_1111100;
		Dminus[720] = 14'b1111111_1111100;
		Dminus[721] = 14'b1111111_1111100;
		Dminus[722] = 14'b1111111_1111100;
		Dminus[723] = 14'b1111111_1111100;
		Dminus[724] = 14'b1111111_1111100;
		Dminus[725] = 14'b1111111_1111100;
		Dminus[726] = 14'b1111111_1111100;
		Dminus[727] = 14'b1111111_1111100;
		Dminus[728] = 14'b1111111_1111100;
		Dminus[729] = 14'b1111111_1111100;
		Dminus[730] = 14'b1111111_1111100;
		Dminus[731] = 14'b1111111_1111100;
		Dminus[732] = 14'b1111111_1111100;
		Dminus[733] = 14'b1111111_1111100;
		Dminus[734] = 14'b1111111_1111100;
		Dminus[735] = 14'b1111111_1111101;
		Dminus[736] = 14'b1111111_1111101;
		Dminus[737] = 14'b1111111_1111101;
		Dminus[738] = 14'b1111111_1111101;
		Dminus[739] = 14'b1111111_1111101;
		Dminus[740] = 14'b1111111_1111101;
		Dminus[741] = 14'b1111111_1111101;
		Dminus[742] = 14'b1111111_1111101;
		Dminus[743] = 14'b1111111_1111101;
		Dminus[744] = 14'b1111111_1111101;
		Dminus[745] = 14'b1111111_1111101;
		Dminus[746] = 14'b1111111_1111101;
		Dminus[747] = 14'b1111111_1111101;
		Dminus[748] = 14'b1111111_1111101;
		Dminus[749] = 14'b1111111_1111101;
		Dminus[750] = 14'b1111111_1111101;
		Dminus[751] = 14'b1111111_1111101;
		Dminus[752] = 14'b1111111_1111101;
		Dminus[753] = 14'b1111111_1111101;
		Dminus[754] = 14'b1111111_1111101;
		Dminus[755] = 14'b1111111_1111101;
		Dminus[756] = 14'b1111111_1111101;
		Dminus[757] = 14'b1111111_1111101;
		Dminus[758] = 14'b1111111_1111101;
		Dminus[759] = 14'b1111111_1111101;
		Dminus[760] = 14'b1111111_1111101;
		Dminus[761] = 14'b1111111_1111101;
		Dminus[762] = 14'b1111111_1111101;
		Dminus[763] = 14'b1111111_1111101;
		Dminus[764] = 14'b1111111_1111101;
		Dminus[765] = 14'b1111111_1111101;
		Dminus[766] = 14'b1111111_1111101;
		Dminus[767] = 14'b1111111_1111101;
		Dminus[768] = 14'b1111111_1111101;
		Dminus[769] = 14'b1111111_1111101;
		Dminus[770] = 14'b1111111_1111101;
		Dminus[771] = 14'b1111111_1111101;
		Dminus[772] = 14'b1111111_1111101;
		Dminus[773] = 14'b1111111_1111101;
		Dminus[774] = 14'b1111111_1111101;
		Dminus[775] = 14'b1111111_1111101;
		Dminus[776] = 14'b1111111_1111101;
		Dminus[777] = 14'b1111111_1111101;
		Dminus[778] = 14'b1111111_1111101;
		Dminus[779] = 14'b1111111_1111101;
		Dminus[780] = 14'b1111111_1111101;
		Dminus[781] = 14'b1111111_1111101;
		Dminus[782] = 14'b1111111_1111101;
		Dminus[783] = 14'b1111111_1111101;
		Dminus[784] = 14'b1111111_1111101;
		Dminus[785] = 14'b1111111_1111101;
		Dminus[786] = 14'b1111111_1111101;
		Dminus[787] = 14'b1111111_1111101;
		Dminus[788] = 14'b1111111_1111101;
		Dminus[789] = 14'b1111111_1111101;
		Dminus[790] = 14'b1111111_1111101;
		Dminus[791] = 14'b1111111_1111101;
		Dminus[792] = 14'b1111111_1111101;
		Dminus[793] = 14'b1111111_1111101;
		Dminus[794] = 14'b1111111_1111101;
		Dminus[795] = 14'b1111111_1111101;
		Dminus[796] = 14'b1111111_1111110;
		Dminus[797] = 14'b1111111_1111110;
		Dminus[798] = 14'b1111111_1111110;
		Dminus[799] = 14'b1111111_1111110;
		Dminus[800] = 14'b1111111_1111110;
		Dminus[801] = 14'b1111111_1111110;
		Dminus[802] = 14'b1111111_1111110;
		Dminus[803] = 14'b1111111_1111110;
		Dminus[804] = 14'b1111111_1111110;
		Dminus[805] = 14'b1111111_1111110;
		Dminus[806] = 14'b1111111_1111110;
		Dminus[807] = 14'b1111111_1111110;
		Dminus[808] = 14'b1111111_1111110;
		Dminus[809] = 14'b1111111_1111110;
		Dminus[810] = 14'b1111111_1111110;
		Dminus[811] = 14'b1111111_1111110;
		Dminus[812] = 14'b1111111_1111110;
		Dminus[813] = 14'b1111111_1111110;
		Dminus[814] = 14'b1111111_1111110;
		Dminus[815] = 14'b1111111_1111110;
		Dminus[816] = 14'b1111111_1111110;
		Dminus[817] = 14'b1111111_1111110;
		Dminus[818] = 14'b1111111_1111110;
		Dminus[819] = 14'b1111111_1111110;
		Dminus[820] = 14'b1111111_1111110;
		Dminus[821] = 14'b1111111_1111110;
		Dminus[822] = 14'b1111111_1111110;
		Dminus[823] = 14'b1111111_1111110;
		Dminus[824] = 14'b1111111_1111110;
		Dminus[825] = 14'b1111111_1111110;
		Dminus[826] = 14'b1111111_1111110;
		Dminus[827] = 14'b1111111_1111110;
		Dminus[828] = 14'b1111111_1111110;
		Dminus[829] = 14'b1111111_1111110;
		Dminus[830] = 14'b1111111_1111110;
		Dminus[831] = 14'b1111111_1111110;
		Dminus[832] = 14'b1111111_1111110;
		Dminus[833] = 14'b1111111_1111110;
		Dminus[834] = 14'b1111111_1111110;
		Dminus[835] = 14'b1111111_1111110;
		Dminus[836] = 14'b1111111_1111110;
		Dminus[837] = 14'b1111111_1111110;
		Dminus[838] = 14'b1111111_1111110;
		Dminus[839] = 14'b1111111_1111110;
		Dminus[840] = 14'b1111111_1111110;
		Dminus[841] = 14'b1111111_1111110;
		Dminus[842] = 14'b1111111_1111110;
		Dminus[843] = 14'b1111111_1111110;
		Dminus[844] = 14'b1111111_1111110;
		Dminus[845] = 14'b1111111_1111110;
		Dminus[846] = 14'b1111111_1111110;
		Dminus[847] = 14'b1111111_1111110;
		Dminus[848] = 14'b1111111_1111110;
		Dminus[849] = 14'b1111111_1111110;
		Dminus[850] = 14'b1111111_1111110;
		Dminus[851] = 14'b1111111_1111110;
		Dminus[852] = 14'b1111111_1111110;
		Dminus[853] = 14'b1111111_1111110;
		Dminus[854] = 14'b1111111_1111110;
		Dminus[855] = 14'b1111111_1111110;
		Dminus[856] = 14'b1111111_1111110;
		Dminus[857] = 14'b1111111_1111110;
		Dminus[858] = 14'b1111111_1111110;
		Dminus[859] = 14'b1111111_1111110;
		Dminus[860] = 14'b1111111_1111110;
		Dminus[861] = 14'b1111111_1111110;
		Dminus[862] = 14'b1111111_1111110;
		Dminus[863] = 14'b1111111_1111110;
		Dminus[864] = 14'b1111111_1111110;
		Dminus[865] = 14'b1111111_1111110;
		Dminus[866] = 14'b1111111_1111110;
		Dminus[867] = 14'b1111111_1111110;
		Dminus[868] = 14'b1111111_1111110;
		Dminus[869] = 14'b1111111_1111110;
		Dminus[870] = 14'b1111111_1111110;
		Dminus[871] = 14'b1111111_1111110;
		Dminus[872] = 14'b1111111_1111110;
		Dminus[873] = 14'b1111111_1111110;
		Dminus[874] = 14'b1111111_1111110;
		Dminus[875] = 14'b1111111_1111110;
		Dminus[876] = 14'b1111111_1111110;
		Dminus[877] = 14'b1111111_1111110;
		Dminus[878] = 14'b1111111_1111110;
		Dminus[879] = 14'b1111111_1111110;
		Dminus[880] = 14'b1111111_1111110;
		Dminus[881] = 14'b1111111_1111110;
		Dminus[882] = 14'b1111111_1111110;
		Dminus[883] = 14'b1111111_1111110;
		Dminus[884] = 14'b1111111_1111110;
		Dminus[885] = 14'b1111111_1111110;
		Dminus[886] = 14'b1111111_1111110;
		Dminus[887] = 14'b1111111_1111110;
		Dminus[888] = 14'b1111111_1111110;
		Dminus[889] = 14'b1111111_1111110;
		Dminus[890] = 14'b1111111_1111111;
		Dminus[891] = 14'b1111111_1111111;
		Dminus[892] = 14'b1111111_1111111;
		Dminus[893] = 14'b1111111_1111111;
		Dminus[894] = 14'b1111111_1111111;
		Dminus[895] = 14'b1111111_1111111;
		Dminus[896] = 14'b1111111_1111111;
		Dminus[897] = 14'b1111111_1111111;
		Dminus[898] = 14'b1111111_1111111;
		Dminus[899] = 14'b1111111_1111111;
		Dminus[900] = 14'b1111111_1111111;
		Dminus[901] = 14'b1111111_1111111;
		Dminus[902] = 14'b1111111_1111111;
		Dminus[903] = 14'b1111111_1111111;
		Dminus[904] = 14'b1111111_1111111;
		Dminus[905] = 14'b1111111_1111111;
		Dminus[906] = 14'b1111111_1111111;
		Dminus[907] = 14'b1111111_1111111;
		Dminus[908] = 14'b1111111_1111111;
		Dminus[909] = 14'b1111111_1111111;
		Dminus[910] = 14'b1111111_1111111;
		Dminus[911] = 14'b1111111_1111111;
		Dminus[912] = 14'b1111111_1111111;
		Dminus[913] = 14'b1111111_1111111;
		Dminus[914] = 14'b1111111_1111111;
		Dminus[915] = 14'b1111111_1111111;
		Dminus[916] = 14'b1111111_1111111;
		Dminus[917] = 14'b1111111_1111111;
		Dminus[918] = 14'b1111111_1111111;
		Dminus[919] = 14'b1111111_1111111;
		Dminus[920] = 14'b1111111_1111111;
		Dminus[921] = 14'b1111111_1111111;
		Dminus[922] = 14'b1111111_1111111;
		Dminus[923] = 14'b1111111_1111111;
		Dminus[924] = 14'b1111111_1111111;
		Dminus[925] = 14'b1111111_1111111;
		Dminus[926] = 14'b1111111_1111111;
		Dminus[927] = 14'b1111111_1111111;
		Dminus[928] = 14'b1111111_1111111;
		Dminus[929] = 14'b1111111_1111111;
		Dminus[930] = 14'b1111111_1111111;
		Dminus[931] = 14'b1111111_1111111;
		Dminus[932] = 14'b1111111_1111111;
		Dminus[933] = 14'b1111111_1111111;
		Dminus[934] = 14'b1111111_1111111;
		Dminus[935] = 14'b1111111_1111111;
		Dminus[936] = 14'b1111111_1111111;
		Dminus[937] = 14'b1111111_1111111;
		Dminus[938] = 14'b1111111_1111111;
		Dminus[939] = 14'b1111111_1111111;
		Dminus[940] = 14'b1111111_1111111;
		Dminus[941] = 14'b1111111_1111111;
		Dminus[942] = 14'b1111111_1111111;
		Dminus[943] = 14'b1111111_1111111;
		Dminus[944] = 14'b1111111_1111111;
		Dminus[945] = 14'b1111111_1111111;
		Dminus[946] = 14'b1111111_1111111;
		Dminus[947] = 14'b1111111_1111111;
		Dminus[948] = 14'b1111111_1111111;
		Dminus[949] = 14'b1111111_1111111;
		Dminus[950] = 14'b1111111_1111111;
		Dminus[951] = 14'b1111111_1111111;
		Dminus[952] = 14'b1111111_1111111;
		Dminus[953] = 14'b1111111_1111111;
		Dminus[954] = 14'b1111111_1111111;
		Dminus[955] = 14'b1111111_1111111;
		Dminus[956] = 14'b1111111_1111111;
		Dminus[957] = 14'b1111111_1111111;
		Dminus[958] = 14'b1111111_1111111;
		Dminus[959] = 14'b1111111_1111111;
		Dminus[960] = 14'b1111111_1111111;
		Dminus[961] = 14'b1111111_1111111;
		Dminus[962] = 14'b1111111_1111111;
		Dminus[963] = 14'b1111111_1111111;
		Dminus[964] = 14'b1111111_1111111;
		Dminus[965] = 14'b1111111_1111111;
		Dminus[966] = 14'b1111111_1111111;
		Dminus[967] = 14'b1111111_1111111;
		Dminus[968] = 14'b1111111_1111111;
		Dminus[969] = 14'b1111111_1111111;
		Dminus[970] = 14'b1111111_1111111;
		Dminus[971] = 14'b1111111_1111111;
		Dminus[972] = 14'b1111111_1111111;
		Dminus[973] = 14'b1111111_1111111;
		Dminus[974] = 14'b1111111_1111111;
		Dminus[975] = 14'b1111111_1111111;
		Dminus[976] = 14'b1111111_1111111;
		Dminus[977] = 14'b1111111_1111111;
		Dminus[978] = 14'b1111111_1111111;
		Dminus[979] = 14'b1111111_1111111;
		Dminus[980] = 14'b1111111_1111111;
		Dminus[981] = 14'b1111111_1111111;
		Dminus[982] = 14'b1111111_1111111;
		Dminus[983] = 14'b1111111_1111111;
		Dminus[984] = 14'b1111111_1111111;
		Dminus[985] = 14'b1111111_1111111;
		Dminus[986] = 14'b1111111_1111111;
		Dminus[987] = 14'b1111111_1111111;
		Dminus[988] = 14'b1111111_1111111;
		Dminus[989] = 14'b1111111_1111111;
		Dminus[990] = 14'b1111111_1111111;
		Dminus[991] = 14'b1111111_1111111;
		Dminus[992] = 14'b1111111_1111111;
		Dminus[993] = 14'b1111111_1111111;
		Dminus[994] = 14'b1111111_1111111;
		Dminus[995] = 14'b1111111_1111111;
		Dminus[996] = 14'b1111111_1111111;
		Dminus[997] = 14'b1111111_1111111;
		Dminus[998] = 14'b1111111_1111111;
		Dminus[999] = 14'b1111111_1111111;
		Dminus[1000] = 14'b1111111_1111111;
		Dminus[1001] = 14'b1111111_1111111;
		Dminus[1002] = 14'b1111111_1111111;
		Dminus[1003] = 14'b1111111_1111111;
		Dminus[1004] = 14'b1111111_1111111;
		Dminus[1005] = 14'b1111111_1111111;
		Dminus[1006] = 14'b1111111_1111111;
		Dminus[1007] = 14'b1111111_1111111;
		Dminus[1008] = 14'b1111111_1111111;
		Dminus[1009] = 14'b1111111_1111111;
		Dminus[1010] = 14'b1111111_1111111;
		Dminus[1011] = 14'b1111111_1111111;
		Dminus[1012] = 14'b1111111_1111111;
		Dminus[1013] = 14'b1111111_1111111;
		Dminus[1014] = 14'b1111111_1111111;
		Dminus[1015] = 14'b1111111_1111111;
		Dminus[1016] = 14'b1111111_1111111;
		Dminus[1017] = 14'b1111111_1111111;
		Dminus[1018] = 14'b1111111_1111111;
		Dminus[1019] = 14'b1111111_1111111;
		Dminus[1020] = 14'b1111111_1111111;
		Dminus[1021] = 14'b1111111_1111111;
		Dminus[1022] = 14'b1111111_1111111;
		Dminus[1023] = 14'b1111111_1111111;
		Dminus[1024] = 14'b1111111_1111111;
		Dminus[1025] = 14'b1111111_1111111;
		Dminus[1026] = 14'b1111111_1111111;
		Dminus[1027] = 14'b1111111_1111111;
		Dminus[1028] = 14'b1111111_1111111;
		Dminus[1029] = 14'b1111111_1111111;
		Dminus[1030] = 14'b1111111_1111111;
		Dminus[1031] = 14'b1111111_1111111;
		Dminus[1032] = 14'b1111111_1111111;
		Dminus[1033] = 14'b1111111_1111111;
		Dminus[1034] = 14'b1111111_1111111;
		Dminus[1035] = 14'b1111111_1111111;
		Dminus[1036] = 14'b1111111_1111111;
		Dminus[1037] = 14'b1111111_1111111;
		Dminus[1038] = 14'b1111111_1111111;
		Dminus[1039] = 14'b1111111_1111111;
		Dminus[1040] = 14'b1111111_1111111;
		Dminus[1041] = 14'b1111111_1111111;
		Dminus[1042] = 14'b1111111_1111111;
		Dminus[1043] = 14'b1111111_1111111;
		Dminus[1044] = 14'b1111111_1111111;
		Dminus[1045] = 14'b1111111_1111111;
		Dminus[1046] = 14'b1111111_1111111;
		Dminus[1047] = 14'b1111111_1111111;
		Dminus[1048] = 14'b1111111_1111111;
		Dminus[1049] = 14'b1111111_1111111;
		Dminus[1050] = 14'b1111111_1111111;
		Dminus[1051] = 14'b1111111_1111111;
		Dminus[1052] = 14'b1111111_1111111;
		Dminus[1053] = 14'b1111111_1111111;
		Dminus[1054] = 14'b1111111_1111111;
		Dminus[1055] = 14'b1111111_1111111;
		Dminus[1056] = 14'b1111111_1111111;
		Dminus[1057] = 14'b1111111_1111111;
		Dminus[1058] = 14'b1111111_1111111;
		Dminus[1059] = 14'b1111111_1111111;
		Dminus[1060] = 14'b1111111_1111111;
		Dminus[1061] = 14'b1111111_1111111;
		Dminus[1062] = 14'b1111111_1111111;
		Dminus[1063] = 14'b1111111_1111111;
		Dminus[1064] = 14'b1111111_1111111;
		Dminus[1065] = 14'b1111111_1111111;
		Dminus[1066] = 14'b1111111_1111111;
		Dminus[1067] = 14'b1111111_1111111;
		Dminus[1068] = 14'b1111111_1111111;
		Dminus[1069] = 14'b1111111_1111111;
		Dminus[1070] = 14'b1111111_1111111;
		Dminus[1071] = 14'b1111111_1111111;
		Dminus[1072] = 14'b1111111_1111111;
		Dminus[1073] = 14'b1111111_1111111;
		Dminus[1074] = 14'b1111111_1111111;
		Dminus[1075] = 14'b1111111_1111111;
		Dminus[1076] = 14'b1111111_1111111;
		Dminus[1077] = 14'b1111111_1111111;
		Dminus[1078] = 14'b1111111_1111111;
		Dminus[1079] = 14'b1111111_1111111;
		Dminus[1080] = 14'b1111111_1111111;
		Dminus[1081] = 14'b1111111_1111111;
		Dminus[1082] = 14'b1111111_1111111;
		Dminus[1083] = 14'b1111111_1111111;
		Dminus[1084] = 14'b1111111_1111111;
		Dminus[1085] = 14'b1111111_1111111;
		Dminus[1086] = 14'b1111111_1111111;
		Dminus[1087] = 14'b1111111_1111111;
		Dminus[1088] = 14'b1111111_1111111;
		Dminus[1089] = 14'b1111111_1111111;
		Dminus[1090] = 14'b1111111_1111111;
		Dminus[1091] = 14'b1111111_1111111;
		Dminus[1092] = 14'b0000000_0000000;
		Dminus[1093] = 14'b0000000_0000000;
		Dminus[1094] = 14'b0000000_0000000;
		Dminus[1095] = 14'b0000000_0000000;
		Dminus[1096] = 14'b0000000_0000000;
		Dminus[1097] = 14'b0000000_0000000;
		Dminus[1098] = 14'b0000000_0000000;
		Dminus[1099] = 14'b0000000_0000000;
		Dminus[1100] = 14'b0000000_0000000;
		Dminus[1101] = 14'b0000000_0000000;
		Dminus[1102] = 14'b0000000_0000000;
		Dminus[1103] = 14'b0000000_0000000;
		Dminus[1104] = 14'b0000000_0000000;
		Dminus[1105] = 14'b0000000_0000000;
		Dminus[1106] = 14'b0000000_0000000;
		Dminus[1107] = 14'b0000000_0000000;
		Dminus[1108] = 14'b0000000_0000000;
		Dminus[1109] = 14'b0000000_0000000;
		Dminus[1110] = 14'b0000000_0000000;
		Dminus[1111] = 14'b0000000_0000000;
		Dminus[1112] = 14'b0000000_0000000;
		Dminus[1113] = 14'b0000000_0000000;
		Dminus[1114] = 14'b0000000_0000000;
		Dminus[1115] = 14'b0000000_0000000;
		Dminus[1116] = 14'b0000000_0000000;
		Dminus[1117] = 14'b0000000_0000000;
		Dminus[1118] = 14'b0000000_0000000;
		Dminus[1119] = 14'b0000000_0000000;
		Dminus[1120] = 14'b0000000_0000000;
		Dminus[1121] = 14'b0000000_0000000;
		Dminus[1122] = 14'b0000000_0000000;
		Dminus[1123] = 14'b0000000_0000000;
		Dminus[1124] = 14'b0000000_0000000;
		Dminus[1125] = 14'b0000000_0000000;
		Dminus[1126] = 14'b0000000_0000000;
		Dminus[1127] = 14'b0000000_0000000;
		Dminus[1128] = 14'b0000000_0000000;
		Dminus[1129] = 14'b0000000_0000000;
		Dminus[1130] = 14'b0000000_0000000;
		Dminus[1131] = 14'b0000000_0000000;
		Dminus[1132] = 14'b0000000_0000000;
		Dminus[1133] = 14'b0000000_0000000;
		Dminus[1134] = 14'b0000000_0000000;
		Dminus[1135] = 14'b0000000_0000000;
		Dminus[1136] = 14'b0000000_0000000;
		Dminus[1137] = 14'b0000000_0000000;
		Dminus[1138] = 14'b0000000_0000000;
		Dminus[1139] = 14'b0000000_0000000;
		Dminus[1140] = 14'b0000000_0000000;
		Dminus[1141] = 14'b0000000_0000000;
		Dminus[1142] = 14'b0000000_0000000;
		Dminus[1143] = 14'b0000000_0000000;
		Dminus[1144] = 14'b0000000_0000000;
		Dminus[1145] = 14'b0000000_0000000;
		Dminus[1146] = 14'b0000000_0000000;
		Dminus[1147] = 14'b0000000_0000000;
		Dminus[1148] = 14'b0000000_0000000;
		Dminus[1149] = 14'b0000000_0000000;
		Dminus[1150] = 14'b0000000_0000000;
		Dminus[1151] = 14'b0000000_0000000;
		Dminus[1152] = 14'b0000000_0000000;
		Dminus[1153] = 14'b0000000_0000000;
		Dminus[1154] = 14'b0000000_0000000;
		Dminus[1155] = 14'b0000000_0000000;
		Dminus[1156] = 14'b0000000_0000000;
		Dminus[1157] = 14'b0000000_0000000;
		Dminus[1158] = 14'b0000000_0000000;
		Dminus[1159] = 14'b0000000_0000000;
		Dminus[1160] = 14'b0000000_0000000;
		Dminus[1161] = 14'b0000000_0000000;
		Dminus[1162] = 14'b0000000_0000000;
		Dminus[1163] = 14'b0000000_0000000;
		Dminus[1164] = 14'b0000000_0000000;
		Dminus[1165] = 14'b0000000_0000000;
		Dminus[1166] = 14'b0000000_0000000;
		Dminus[1167] = 14'b0000000_0000000;
		Dminus[1168] = 14'b0000000_0000000;
		Dminus[1169] = 14'b0000000_0000000;
		Dminus[1170] = 14'b0000000_0000000;
		Dminus[1171] = 14'b0000000_0000000;
		Dminus[1172] = 14'b0000000_0000000;
		Dminus[1173] = 14'b0000000_0000000;
		Dminus[1174] = 14'b0000000_0000000;
		Dminus[1175] = 14'b0000000_0000000;
		Dminus[1176] = 14'b0000000_0000000;
		Dminus[1177] = 14'b0000000_0000000;
		Dminus[1178] = 14'b0000000_0000000;
		Dminus[1179] = 14'b0000000_0000000;
		Dminus[1180] = 14'b0000000_0000000;
		Dminus[1181] = 14'b0000000_0000000;
		Dminus[1182] = 14'b0000000_0000000;
		Dminus[1183] = 14'b0000000_0000000;
		Dminus[1184] = 14'b0000000_0000000;
		Dminus[1185] = 14'b0000000_0000000;
		Dminus[1186] = 14'b0000000_0000000;
		Dminus[1187] = 14'b0000000_0000000;
		Dminus[1188] = 14'b0000000_0000000;
		Dminus[1189] = 14'b0000000_0000000;
		Dminus[1190] = 14'b0000000_0000000;
		Dminus[1191] = 14'b0000000_0000000;
		Dminus[1192] = 14'b0000000_0000000;
		Dminus[1193] = 14'b0000000_0000000;
		Dminus[1194] = 14'b0000000_0000000;
		Dminus[1195] = 14'b0000000_0000000;
		Dminus[1196] = 14'b0000000_0000000;
		Dminus[1197] = 14'b0000000_0000000;
		Dminus[1198] = 14'b0000000_0000000;
		Dminus[1199] = 14'b0000000_0000000;
		Dminus[1200] = 14'b0000000_0000000;
		Dminus[1201] = 14'b0000000_0000000;
		Dminus[1202] = 14'b0000000_0000000;
		Dminus[1203] = 14'b0000000_0000000;
		Dminus[1204] = 14'b0000000_0000000;
		Dminus[1205] = 14'b0000000_0000000;
		Dminus[1206] = 14'b0000000_0000000;
		Dminus[1207] = 14'b0000000_0000000;
		Dminus[1208] = 14'b0000000_0000000;
		Dminus[1209] = 14'b0000000_0000000;
		Dminus[1210] = 14'b0000000_0000000;
		Dminus[1211] = 14'b0000000_0000000;
		Dminus[1212] = 14'b0000000_0000000;
		Dminus[1213] = 14'b0000000_0000000;
		Dminus[1214] = 14'b0000000_0000000;
		Dminus[1215] = 14'b0000000_0000000;
		Dminus[1216] = 14'b0000000_0000000;
		Dminus[1217] = 14'b0000000_0000000;
		Dminus[1218] = 14'b0000000_0000000;
		Dminus[1219] = 14'b0000000_0000000;
		Dminus[1220] = 14'b0000000_0000000;
		Dminus[1221] = 14'b0000000_0000000;
		Dminus[1222] = 14'b0000000_0000000;
		Dminus[1223] = 14'b0000000_0000000;
		Dminus[1224] = 14'b0000000_0000000;
		Dminus[1225] = 14'b0000000_0000000;
		Dminus[1226] = 14'b0000000_0000000;
		Dminus[1227] = 14'b0000000_0000000;
		Dminus[1228] = 14'b0000000_0000000;
		Dminus[1229] = 14'b0000000_0000000;
		Dminus[1230] = 14'b0000000_0000000;
		Dminus[1231] = 14'b0000000_0000000;
		Dminus[1232] = 14'b0000000_0000000;
		Dminus[1233] = 14'b0000000_0000000;
		Dminus[1234] = 14'b0000000_0000000;
		Dminus[1235] = 14'b0000000_0000000;
		Dminus[1236] = 14'b0000000_0000000;
		Dminus[1237] = 14'b0000000_0000000;
		Dminus[1238] = 14'b0000000_0000000;
		Dminus[1239] = 14'b0000000_0000000;
		Dminus[1240] = 14'b0000000_0000000;
		Dminus[1241] = 14'b0000000_0000000;
		Dminus[1242] = 14'b0000000_0000000;
		Dminus[1243] = 14'b0000000_0000000;
		Dminus[1244] = 14'b0000000_0000000;
		Dminus[1245] = 14'b0000000_0000000;
		Dminus[1246] = 14'b0000000_0000000;
		Dminus[1247] = 14'b0000000_0000000;
		Dminus[1248] = 14'b0000000_0000000;
		Dminus[1249] = 14'b0000000_0000000;
		Dminus[1250] = 14'b0000000_0000000;
		Dminus[1251] = 14'b0000000_0000000;
		Dminus[1252] = 14'b0000000_0000000;
		Dminus[1253] = 14'b0000000_0000000;
		Dminus[1254] = 14'b0000000_0000000;
		Dminus[1255] = 14'b0000000_0000000;
		Dminus[1256] = 14'b0000000_0000000;
		Dminus[1257] = 14'b0000000_0000000;
		Dminus[1258] = 14'b0000000_0000000;
		Dminus[1259] = 14'b0000000_0000000;
		Dminus[1260] = 14'b0000000_0000000;
		Dminus[1261] = 14'b0000000_0000000;
		Dminus[1262] = 14'b0000000_0000000;
		Dminus[1263] = 14'b0000000_0000000;
		Dminus[1264] = 14'b0000000_0000000;
		Dminus[1265] = 14'b0000000_0000000;
		Dminus[1266] = 14'b0000000_0000000;
		Dminus[1267] = 14'b0000000_0000000;
		Dminus[1268] = 14'b0000000_0000000;
		Dminus[1269] = 14'b0000000_0000000;
		Dminus[1270] = 14'b0000000_0000000;
		Dminus[1271] = 14'b0000000_0000000;
		Dminus[1272] = 14'b0000000_0000000;
		Dminus[1273] = 14'b0000000_0000000;
		Dminus[1274] = 14'b0000000_0000000;
		Dminus[1275] = 14'b0000000_0000000;
		Dminus[1276] = 14'b0000000_0000000;
		Dminus[1277] = 14'b0000000_0000000;
		Dminus[1278] = 14'b0000000_0000000;
		Dminus[1279] = 14'b0000000_0000000;
		Dminus[1280] = 14'b0000000_0000000;
		Dminus[1281] = 14'b0000000_0000000;
		Dminus[1282] = 14'b0000000_0000000;
		Dminus[1283] = 14'b0000000_0000000;
		Dminus[1284] = 14'b0000000_0000000;
		Dminus[1285] = 14'b0000000_0000000;
		Dminus[1286] = 14'b0000000_0000000;
		Dminus[1287] = 14'b0000000_0000000;
		Dminus[1288] = 14'b0000000_0000000;
		Dminus[1289] = 14'b0000000_0000000;
		Dminus[1290] = 14'b0000000_0000000;
		Dminus[1291] = 14'b0000000_0000000;
		Dminus[1292] = 14'b0000000_0000000;
		Dminus[1293] = 14'b0000000_0000000;
		Dminus[1294] = 14'b0000000_0000000;
		Dminus[1295] = 14'b0000000_0000000;
		Dminus[1296] = 14'b0000000_0000000;
		Dminus[1297] = 14'b0000000_0000000;
		Dminus[1298] = 14'b0000000_0000000;
		Dminus[1299] = 14'b0000000_0000000;
		Dminus[1300] = 14'b0000000_0000000;
		Dminus[1301] = 14'b0000000_0000000;
		Dminus[1302] = 14'b0000000_0000000;
		Dminus[1303] = 14'b0000000_0000000;
		Dminus[1304] = 14'b0000000_0000000;
		Dminus[1305] = 14'b0000000_0000000;
		Dminus[1306] = 14'b0000000_0000000;
		Dminus[1307] = 14'b0000000_0000000;
		Dminus[1308] = 14'b0000000_0000000;
		Dminus[1309] = 14'b0000000_0000000;
		Dminus[1310] = 14'b0000000_0000000;
		Dminus[1311] = 14'b0000000_0000000;
		Dminus[1312] = 14'b0000000_0000000;
		Dminus[1313] = 14'b0000000_0000000;
		Dminus[1314] = 14'b0000000_0000000;
		Dminus[1315] = 14'b0000000_0000000;
		Dminus[1316] = 14'b0000000_0000000;
		Dminus[1317] = 14'b0000000_0000000;
		Dminus[1318] = 14'b0000000_0000000;
		Dminus[1319] = 14'b0000000_0000000;
		Dminus[1320] = 14'b0000000_0000000;
		Dminus[1321] = 14'b0000000_0000000;
		Dminus[1322] = 14'b0000000_0000000;
		Dminus[1323] = 14'b0000000_0000000;
		Dminus[1324] = 14'b0000000_0000000;
		Dminus[1325] = 14'b0000000_0000000;
		Dminus[1326] = 14'b0000000_0000000;
		Dminus[1327] = 14'b0000000_0000000;
		Dminus[1328] = 14'b0000000_0000000;
		Dminus[1329] = 14'b0000000_0000000;
		Dminus[1330] = 14'b0000000_0000000;
		Dminus[1331] = 14'b0000000_0000000;
		Dminus[1332] = 14'b0000000_0000000;
		Dminus[1333] = 14'b0000000_0000000;
		Dminus[1334] = 14'b0000000_0000000;
		Dminus[1335] = 14'b0000000_0000000;
		Dminus[1336] = 14'b0000000_0000000;
		Dminus[1337] = 14'b0000000_0000000;
		Dminus[1338] = 14'b0000000_0000000;
		Dminus[1339] = 14'b0000000_0000000;
		Dminus[1340] = 14'b0000000_0000000;
		Dminus[1341] = 14'b0000000_0000000;
		Dminus[1342] = 14'b0000000_0000000;
		Dminus[1343] = 14'b0000000_0000000;
		Dminus[1344] = 14'b0000000_0000000;
		Dminus[1345] = 14'b0000000_0000000;
		Dminus[1346] = 14'b0000000_0000000;
		Dminus[1347] = 14'b0000000_0000000;
		Dminus[1348] = 14'b0000000_0000000;
		Dminus[1349] = 14'b0000000_0000000;
		Dminus[1350] = 14'b0000000_0000000;
		Dminus[1351] = 14'b0000000_0000000;
		Dminus[1352] = 14'b0000000_0000000;
		Dminus[1353] = 14'b0000000_0000000;
		Dminus[1354] = 14'b0000000_0000000;
		Dminus[1355] = 14'b0000000_0000000;
		Dminus[1356] = 14'b0000000_0000000;
		Dminus[1357] = 14'b0000000_0000000;
		Dminus[1358] = 14'b0000000_0000000;
		Dminus[1359] = 14'b0000000_0000000;
		Dminus[1360] = 14'b0000000_0000000;
		Dminus[1361] = 14'b0000000_0000000;
		Dminus[1362] = 14'b0000000_0000000;
		Dminus[1363] = 14'b0000000_0000000;
		Dminus[1364] = 14'b0000000_0000000;
		Dminus[1365] = 14'b0000000_0000000;
		Dminus[1366] = 14'b0000000_0000000;
		Dminus[1367] = 14'b0000000_0000000;
		Dminus[1368] = 14'b0000000_0000000;
		Dminus[1369] = 14'b0000000_0000000;
		Dminus[1370] = 14'b0000000_0000000;
		Dminus[1371] = 14'b0000000_0000000;
		Dminus[1372] = 14'b0000000_0000000;
		Dminus[1373] = 14'b0000000_0000000;
		Dminus[1374] = 14'b0000000_0000000;
		Dminus[1375] = 14'b0000000_0000000;
		Dminus[1376] = 14'b0000000_0000000;
		Dminus[1377] = 14'b0000000_0000000;
		Dminus[1378] = 14'b0000000_0000000;
		Dminus[1379] = 14'b0000000_0000000;
		Dminus[1380] = 14'b0000000_0000000;
		Dminus[1381] = 14'b0000000_0000000;
		Dminus[1382] = 14'b0000000_0000000;
		Dminus[1383] = 14'b0000000_0000000;
		Dminus[1384] = 14'b0000000_0000000;
		Dminus[1385] = 14'b0000000_0000000;
		Dminus[1386] = 14'b0000000_0000000;
		Dminus[1387] = 14'b0000000_0000000;
		Dminus[1388] = 14'b0000000_0000000;
		Dminus[1389] = 14'b0000000_0000000;
		Dminus[1390] = 14'b0000000_0000000;
		Dminus[1391] = 14'b0000000_0000000;
		Dminus[1392] = 14'b0000000_0000000;
		Dminus[1393] = 14'b0000000_0000000;
		Dminus[1394] = 14'b0000000_0000000;
		Dminus[1395] = 14'b0000000_0000000;
		Dminus[1396] = 14'b0000000_0000000;
		Dminus[1397] = 14'b0000000_0000000;
		Dminus[1398] = 14'b0000000_0000000;
		Dminus[1399] = 14'b0000000_0000000;
		Dminus[1400] = 14'b0000000_0000000;
		Dminus[1401] = 14'b0000000_0000000;
		Dminus[1402] = 14'b0000000_0000000;
		Dminus[1403] = 14'b0000000_0000000;
		Dminus[1404] = 14'b0000000_0000000;
		Dminus[1405] = 14'b0000000_0000000;
		Dminus[1406] = 14'b0000000_0000000;
		Dminus[1407] = 14'b0000000_0000000;
		Dminus[1408] = 14'b0000000_0000000;
		Dminus[1409] = 14'b0000000_0000000;
		Dminus[1410] = 14'b0000000_0000000;
		Dminus[1411] = 14'b0000000_0000000;
		Dminus[1412] = 14'b0000000_0000000;
		Dminus[1413] = 14'b0000000_0000000;
		Dminus[1414] = 14'b0000000_0000000;
		Dminus[1415] = 14'b0000000_0000000;
		Dminus[1416] = 14'b0000000_0000000;
		Dminus[1417] = 14'b0000000_0000000;
		Dminus[1418] = 14'b0000000_0000000;
		Dminus[1419] = 14'b0000000_0000000;
		Dminus[1420] = 14'b0000000_0000000;
		Dminus[1421] = 14'b0000000_0000000;
		Dminus[1422] = 14'b0000000_0000000;
		Dminus[1423] = 14'b0000000_0000000;
		Dminus[1424] = 14'b0000000_0000000;
		Dminus[1425] = 14'b0000000_0000000;
		Dminus[1426] = 14'b0000000_0000000;
		Dminus[1427] = 14'b0000000_0000000;
		Dminus[1428] = 14'b0000000_0000000;
		Dminus[1429] = 14'b0000000_0000000;
		Dminus[1430] = 14'b0000000_0000000;
		Dminus[1431] = 14'b0000000_0000000;
		Dminus[1432] = 14'b0000000_0000000;
		Dminus[1433] = 14'b0000000_0000000;
		Dminus[1434] = 14'b0000000_0000000;
		Dminus[1435] = 14'b0000000_0000000;
		Dminus[1436] = 14'b0000000_0000000;
		Dminus[1437] = 14'b0000000_0000000;
		Dminus[1438] = 14'b0000000_0000000;
		Dminus[1439] = 14'b0000000_0000000;
		Dminus[1440] = 14'b0000000_0000000;
		Dminus[1441] = 14'b0000000_0000000;
		Dminus[1442] = 14'b0000000_0000000;
		Dminus[1443] = 14'b0000000_0000000;
		Dminus[1444] = 14'b0000000_0000000;
		Dminus[1445] = 14'b0000000_0000000;
		Dminus[1446] = 14'b0000000_0000000;
		Dminus[1447] = 14'b0000000_0000000;
		Dminus[1448] = 14'b0000000_0000000;
		Dminus[1449] = 14'b0000000_0000000;
		Dminus[1450] = 14'b0000000_0000000;
		Dminus[1451] = 14'b0000000_0000000;
		Dminus[1452] = 14'b0000000_0000000;
		Dminus[1453] = 14'b0000000_0000000;
		Dminus[1454] = 14'b0000000_0000000;
		Dminus[1455] = 14'b0000000_0000000;
		Dminus[1456] = 14'b0000000_0000000;
		Dminus[1457] = 14'b0000000_0000000;
		Dminus[1458] = 14'b0000000_0000000;
		Dminus[1459] = 14'b0000000_0000000;
		Dminus[1460] = 14'b0000000_0000000;
		Dminus[1461] = 14'b0000000_0000000;
		Dminus[1462] = 14'b0000000_0000000;
		Dminus[1463] = 14'b0000000_0000000;
		Dminus[1464] = 14'b0000000_0000000;
		Dminus[1465] = 14'b0000000_0000000;
		Dminus[1466] = 14'b0000000_0000000;
		Dminus[1467] = 14'b0000000_0000000;
		Dminus[1468] = 14'b0000000_0000000;
		Dminus[1469] = 14'b0000000_0000000;
		Dminus[1470] = 14'b0000000_0000000;
		Dminus[1471] = 14'b0000000_0000000;
		Dminus[1472] = 14'b0000000_0000000;
		Dminus[1473] = 14'b0000000_0000000;
		Dminus[1474] = 14'b0000000_0000000;
		Dminus[1475] = 14'b0000000_0000000;
		Dminus[1476] = 14'b0000000_0000000;
		Dminus[1477] = 14'b0000000_0000000;
		Dminus[1478] = 14'b0000000_0000000;
		Dminus[1479] = 14'b0000000_0000000;
		Dminus[1480] = 14'b0000000_0000000;
		Dminus[1481] = 14'b0000000_0000000;
		Dminus[1482] = 14'b0000000_0000000;
		Dminus[1483] = 14'b0000000_0000000;
		Dminus[1484] = 14'b0000000_0000000;
		Dminus[1485] = 14'b0000000_0000000;
		Dminus[1486] = 14'b0000000_0000000;
		Dminus[1487] = 14'b0000000_0000000;
		Dminus[1488] = 14'b0000000_0000000;
		Dminus[1489] = 14'b0000000_0000000;
		Dminus[1490] = 14'b0000000_0000000;
		Dminus[1491] = 14'b0000000_0000000;
		Dminus[1492] = 14'b0000000_0000000;
		Dminus[1493] = 14'b0000000_0000000;
		Dminus[1494] = 14'b0000000_0000000;
		Dminus[1495] = 14'b0000000_0000000;
		Dminus[1496] = 14'b0000000_0000000;
		Dminus[1497] = 14'b0000000_0000000;
		Dminus[1498] = 14'b0000000_0000000;
		Dminus[1499] = 14'b0000000_0000000;
		Dminus[1500] = 14'b0000000_0000000;
		Dminus[1501] = 14'b0000000_0000000;
		Dminus[1502] = 14'b0000000_0000000;
		Dminus[1503] = 14'b0000000_0000000;
		Dminus[1504] = 14'b0000000_0000000;
		Dminus[1505] = 14'b0000000_0000000;
		Dminus[1506] = 14'b0000000_0000000;
		Dminus[1507] = 14'b0000000_0000000;
		Dminus[1508] = 14'b0000000_0000000;
		Dminus[1509] = 14'b0000000_0000000;
		Dminus[1510] = 14'b0000000_0000000;
		Dminus[1511] = 14'b0000000_0000000;
		Dminus[1512] = 14'b0000000_0000000;
		Dminus[1513] = 14'b0000000_0000000;
		Dminus[1514] = 14'b0000000_0000000;
		Dminus[1515] = 14'b0000000_0000000;
		Dminus[1516] = 14'b0000000_0000000;
		Dminus[1517] = 14'b0000000_0000000;
		Dminus[1518] = 14'b0000000_0000000;
		Dminus[1519] = 14'b0000000_0000000;
		Dminus[1520] = 14'b0000000_0000000;
		Dminus[1521] = 14'b0000000_0000000;
		Dminus[1522] = 14'b0000000_0000000;
		Dminus[1523] = 14'b0000000_0000000;
		Dminus[1524] = 14'b0000000_0000000;
		Dminus[1525] = 14'b0000000_0000000;
		Dminus[1526] = 14'b0000000_0000000;
		Dminus[1527] = 14'b0000000_0000000;
		Dminus[1528] = 14'b0000000_0000000;
		Dminus[1529] = 14'b0000000_0000000;
		Dminus[1530] = 14'b0000000_0000000;
		Dminus[1531] = 14'b0000000_0000000;
		Dminus[1532] = 14'b0000000_0000000;
		Dminus[1533] = 14'b0000000_0000000;
		Dminus[1534] = 14'b0000000_0000000;
		Dminus[1535] = 14'b0000000_0000000;
		Dminus[1536] = 14'b0000000_0000000;
		Dminus[1537] = 14'b0000000_0000000;
		Dminus[1538] = 14'b0000000_0000000;
		Dminus[1539] = 14'b0000000_0000000;
		Dminus[1540] = 14'b0000000_0000000;
		Dminus[1541] = 14'b0000000_0000000;
		Dminus[1542] = 14'b0000000_0000000;
		Dminus[1543] = 14'b0000000_0000000;
		Dminus[1544] = 14'b0000000_0000000;
		Dminus[1545] = 14'b0000000_0000000;
		Dminus[1546] = 14'b0000000_0000000;
		Dminus[1547] = 14'b0000000_0000000;
		Dminus[1548] = 14'b0000000_0000000;
		Dminus[1549] = 14'b0000000_0000000;
		Dminus[1550] = 14'b0000000_0000000;
		Dminus[1551] = 14'b0000000_0000000;
		Dminus[1552] = 14'b0000000_0000000;
		Dminus[1553] = 14'b0000000_0000000;
		Dminus[1554] = 14'b0000000_0000000;
		Dminus[1555] = 14'b0000000_0000000;
		Dminus[1556] = 14'b0000000_0000000;
		Dminus[1557] = 14'b0000000_0000000;
		Dminus[1558] = 14'b0000000_0000000;
		Dminus[1559] = 14'b0000000_0000000;
		Dminus[1560] = 14'b0000000_0000000;
		Dminus[1561] = 14'b0000000_0000000;
		Dminus[1562] = 14'b0000000_0000000;
		Dminus[1563] = 14'b0000000_0000000;
		Dminus[1564] = 14'b0000000_0000000;
		Dminus[1565] = 14'b0000000_0000000;
		Dminus[1566] = 14'b0000000_0000000;
		Dminus[1567] = 14'b0000000_0000000;
		Dminus[1568] = 14'b0000000_0000000;
		Dminus[1569] = 14'b0000000_0000000;
		Dminus[1570] = 14'b0000000_0000000;
		Dminus[1571] = 14'b0000000_0000000;
		Dminus[1572] = 14'b0000000_0000000;
		Dminus[1573] = 14'b0000000_0000000;
		Dminus[1574] = 14'b0000000_0000000;
		Dminus[1575] = 14'b0000000_0000000;
		Dminus[1576] = 14'b0000000_0000000;
		Dminus[1577] = 14'b0000000_0000000;
		Dminus[1578] = 14'b0000000_0000000;
		Dminus[1579] = 14'b0000000_0000000;
		Dminus[1580] = 14'b0000000_0000000;
		Dminus[1581] = 14'b0000000_0000000;
		Dminus[1582] = 14'b0000000_0000000;
		Dminus[1583] = 14'b0000000_0000000;
		Dminus[1584] = 14'b0000000_0000000;
		Dminus[1585] = 14'b0000000_0000000;
		Dminus[1586] = 14'b0000000_0000000;
		Dminus[1587] = 14'b0000000_0000000;
		Dminus[1588] = 14'b0000000_0000000;
		Dminus[1589] = 14'b0000000_0000000;
		Dminus[1590] = 14'b0000000_0000000;
		Dminus[1591] = 14'b0000000_0000000;
		Dminus[1592] = 14'b0000000_0000000;
		Dminus[1593] = 14'b0000000_0000000;
		Dminus[1594] = 14'b0000000_0000000;
		Dminus[1595] = 14'b0000000_0000000;
		Dminus[1596] = 14'b0000000_0000000;
		Dminus[1597] = 14'b0000000_0000000;
		Dminus[1598] = 14'b0000000_0000000;
		Dminus[1599] = 14'b0000000_0000000;
		Dminus[1600] = 14'b0000000_0000000;
		Dminus[1601] = 14'b0000000_0000000;
		Dminus[1602] = 14'b0000000_0000000;
		Dminus[1603] = 14'b0000000_0000000;
		Dminus[1604] = 14'b0000000_0000000;
		Dminus[1605] = 14'b0000000_0000000;
		Dminus[1606] = 14'b0000000_0000000;
		Dminus[1607] = 14'b0000000_0000000;
		Dminus[1608] = 14'b0000000_0000000;
		Dminus[1609] = 14'b0000000_0000000;
		Dminus[1610] = 14'b0000000_0000000;
		Dminus[1611] = 14'b0000000_0000000;
		Dminus[1612] = 14'b0000000_0000000;
		Dminus[1613] = 14'b0000000_0000000;
		Dminus[1614] = 14'b0000000_0000000;
		Dminus[1615] = 14'b0000000_0000000;
		Dminus[1616] = 14'b0000000_0000000;
		Dminus[1617] = 14'b0000000_0000000;
		Dminus[1618] = 14'b0000000_0000000;
		Dminus[1619] = 14'b0000000_0000000;
		Dminus[1620] = 14'b0000000_0000000;
		Dminus[1621] = 14'b0000000_0000000;
		Dminus[1622] = 14'b0000000_0000000;
		Dminus[1623] = 14'b0000000_0000000;
		Dminus[1624] = 14'b0000000_0000000;
		Dminus[1625] = 14'b0000000_0000000;
		Dminus[1626] = 14'b0000000_0000000;
		Dminus[1627] = 14'b0000000_0000000;
		Dminus[1628] = 14'b0000000_0000000;
		Dminus[1629] = 14'b0000000_0000000;
		Dminus[1630] = 14'b0000000_0000000;
		Dminus[1631] = 14'b0000000_0000000;
		Dminus[1632] = 14'b0000000_0000000;
		Dminus[1633] = 14'b0000000_0000000;
		Dminus[1634] = 14'b0000000_0000000;
		Dminus[1635] = 14'b0000000_0000000;
		Dminus[1636] = 14'b0000000_0000000;
		Dminus[1637] = 14'b0000000_0000000;
		Dminus[1638] = 14'b0000000_0000000;
		Dminus[1639] = 14'b0000000_0000000;
		Dminus[1640] = 14'b0000000_0000000;
		Dminus[1641] = 14'b0000000_0000000;
		Dminus[1642] = 14'b0000000_0000000;
		Dminus[1643] = 14'b0000000_0000000;
		Dminus[1644] = 14'b0000000_0000000;
		Dminus[1645] = 14'b0000000_0000000;
		Dminus[1646] = 14'b0000000_0000000;
		Dminus[1647] = 14'b0000000_0000000;
		Dminus[1648] = 14'b0000000_0000000;
		Dminus[1649] = 14'b0000000_0000000;
		Dminus[1650] = 14'b0000000_0000000;
		Dminus[1651] = 14'b0000000_0000000;
		Dminus[1652] = 14'b0000000_0000000;
		Dminus[1653] = 14'b0000000_0000000;
		Dminus[1654] = 14'b0000000_0000000;
		Dminus[1655] = 14'b0000000_0000000;
		Dminus[1656] = 14'b0000000_0000000;
		Dminus[1657] = 14'b0000000_0000000;
		Dminus[1658] = 14'b0000000_0000000;
		Dminus[1659] = 14'b0000000_0000000;
		Dminus[1660] = 14'b0000000_0000000;
		Dminus[1661] = 14'b0000000_0000000;
		Dminus[1662] = 14'b0000000_0000000;
		Dminus[1663] = 14'b0000000_0000000;
		Dminus[1664] = 14'b0000000_0000000;
		Dminus[1665] = 14'b0000000_0000000;
		Dminus[1666] = 14'b0000000_0000000;
		Dminus[1667] = 14'b0000000_0000000;
		Dminus[1668] = 14'b0000000_0000000;
		Dminus[1669] = 14'b0000000_0000000;
		Dminus[1670] = 14'b0000000_0000000;
		Dminus[1671] = 14'b0000000_0000000;
		Dminus[1672] = 14'b0000000_0000000;
		Dminus[1673] = 14'b0000000_0000000;
		Dminus[1674] = 14'b0000000_0000000;
		Dminus[1675] = 14'b0000000_0000000;
		Dminus[1676] = 14'b0000000_0000000;
		Dminus[1677] = 14'b0000000_0000000;
		Dminus[1678] = 14'b0000000_0000000;
		Dminus[1679] = 14'b0000000_0000000;
		Dminus[1680] = 14'b0000000_0000000;
		Dminus[1681] = 14'b0000000_0000000;
		Dminus[1682] = 14'b0000000_0000000;
		Dminus[1683] = 14'b0000000_0000000;
		Dminus[1684] = 14'b0000000_0000000;
		Dminus[1685] = 14'b0000000_0000000;
		Dminus[1686] = 14'b0000000_0000000;
		Dminus[1687] = 14'b0000000_0000000;
		Dminus[1688] = 14'b0000000_0000000;
		Dminus[1689] = 14'b0000000_0000000;
		Dminus[1690] = 14'b0000000_0000000;
		Dminus[1691] = 14'b0000000_0000000;
		Dminus[1692] = 14'b0000000_0000000;
		Dminus[1693] = 14'b0000000_0000000;
		Dminus[1694] = 14'b0000000_0000000;
		Dminus[1695] = 14'b0000000_0000000;
		Dminus[1696] = 14'b0000000_0000000;
		Dminus[1697] = 14'b0000000_0000000;
		Dminus[1698] = 14'b0000000_0000000;
		Dminus[1699] = 14'b0000000_0000000;
		Dminus[1700] = 14'b0000000_0000000;
		Dminus[1701] = 14'b0000000_0000000;
		Dminus[1702] = 14'b0000000_0000000;
		Dminus[1703] = 14'b0000000_0000000;
		Dminus[1704] = 14'b0000000_0000000;
		Dminus[1705] = 14'b0000000_0000000;
		Dminus[1706] = 14'b0000000_0000000;
		Dminus[1707] = 14'b0000000_0000000;
		Dminus[1708] = 14'b0000000_0000000;
		Dminus[1709] = 14'b0000000_0000000;
		Dminus[1710] = 14'b0000000_0000000;
		Dminus[1711] = 14'b0000000_0000000;
		Dminus[1712] = 14'b0000000_0000000;
		Dminus[1713] = 14'b0000000_0000000;
		Dminus[1714] = 14'b0000000_0000000;
		Dminus[1715] = 14'b0000000_0000000;
		Dminus[1716] = 14'b0000000_0000000;
		Dminus[1717] = 14'b0000000_0000000;
		Dminus[1718] = 14'b0000000_0000000;
		Dminus[1719] = 14'b0000000_0000000;
		Dminus[1720] = 14'b0000000_0000000;
		Dminus[1721] = 14'b0000000_0000000;
		Dminus[1722] = 14'b0000000_0000000;
		Dminus[1723] = 14'b0000000_0000000;
		Dminus[1724] = 14'b0000000_0000000;
		Dminus[1725] = 14'b0000000_0000000;
		Dminus[1726] = 14'b0000000_0000000;
		Dminus[1727] = 14'b0000000_0000000;
		Dminus[1728] = 14'b0000000_0000000;
		Dminus[1729] = 14'b0000000_0000000;
		Dminus[1730] = 14'b0000000_0000000;
		Dminus[1731] = 14'b0000000_0000000;
		Dminus[1732] = 14'b0000000_0000000;
		Dminus[1733] = 14'b0000000_0000000;
		Dminus[1734] = 14'b0000000_0000000;
		Dminus[1735] = 14'b0000000_0000000;
		Dminus[1736] = 14'b0000000_0000000;
		Dminus[1737] = 14'b0000000_0000000;
		Dminus[1738] = 14'b0000000_0000000;
		Dminus[1739] = 14'b0000000_0000000;
		Dminus[1740] = 14'b0000000_0000000;
		Dminus[1741] = 14'b0000000_0000000;
		Dminus[1742] = 14'b0000000_0000000;
		Dminus[1743] = 14'b0000000_0000000;
		Dminus[1744] = 14'b0000000_0000000;
		Dminus[1745] = 14'b0000000_0000000;
		Dminus[1746] = 14'b0000000_0000000;
		Dminus[1747] = 14'b0000000_0000000;
		Dminus[1748] = 14'b0000000_0000000;
		Dminus[1749] = 14'b0000000_0000000;
		Dminus[1750] = 14'b0000000_0000000;
		Dminus[1751] = 14'b0000000_0000000;
		Dminus[1752] = 14'b0000000_0000000;
		Dminus[1753] = 14'b0000000_0000000;
		Dminus[1754] = 14'b0000000_0000000;
		Dminus[1755] = 14'b0000000_0000000;
		Dminus[1756] = 14'b0000000_0000000;
		Dminus[1757] = 14'b0000000_0000000;
		Dminus[1758] = 14'b0000000_0000000;
		Dminus[1759] = 14'b0000000_0000000;
		Dminus[1760] = 14'b0000000_0000000;
		Dminus[1761] = 14'b0000000_0000000;
		Dminus[1762] = 14'b0000000_0000000;
		Dminus[1763] = 14'b0000000_0000000;
		Dminus[1764] = 14'b0000000_0000000;
		Dminus[1765] = 14'b0000000_0000000;
		Dminus[1766] = 14'b0000000_0000000;
		Dminus[1767] = 14'b0000000_0000000;
		Dminus[1768] = 14'b0000000_0000000;
		Dminus[1769] = 14'b0000000_0000000;
		Dminus[1770] = 14'b0000000_0000000;
		Dminus[1771] = 14'b0000000_0000000;
		Dminus[1772] = 14'b0000000_0000000;
		Dminus[1773] = 14'b0000000_0000000;
		Dminus[1774] = 14'b0000000_0000000;
		Dminus[1775] = 14'b0000000_0000000;
		Dminus[1776] = 14'b0000000_0000000;
		Dminus[1777] = 14'b0000000_0000000;
		Dminus[1778] = 14'b0000000_0000000;
		Dminus[1779] = 14'b0000000_0000000;
		Dminus[1780] = 14'b0000000_0000000;
		Dminus[1781] = 14'b0000000_0000000;
		Dminus[1782] = 14'b0000000_0000000;
		Dminus[1783] = 14'b0000000_0000000;
		Dminus[1784] = 14'b0000000_0000000;
		Dminus[1785] = 14'b0000000_0000000;
		Dminus[1786] = 14'b0000000_0000000;
		Dminus[1787] = 14'b0000000_0000000;
		Dminus[1788] = 14'b0000000_0000000;
		Dminus[1789] = 14'b0000000_0000000;
		Dminus[1790] = 14'b0000000_0000000;
		Dminus[1791] = 14'b0000000_0000000;
		Dminus[1792] = 14'b0000000_0000000;
		Dminus[1793] = 14'b0000000_0000000;
		Dminus[1794] = 14'b0000000_0000000;
		Dminus[1795] = 14'b0000000_0000000;
		Dminus[1796] = 14'b0000000_0000000;
		Dminus[1797] = 14'b0000000_0000000;
		Dminus[1798] = 14'b0000000_0000000;
		Dminus[1799] = 14'b0000000_0000000;
		Dminus[1800] = 14'b0000000_0000000;
		Dminus[1801] = 14'b0000000_0000000;
		Dminus[1802] = 14'b0000000_0000000;
		Dminus[1803] = 14'b0000000_0000000;
		Dminus[1804] = 14'b0000000_0000000;
		Dminus[1805] = 14'b0000000_0000000;
		Dminus[1806] = 14'b0000000_0000000;
		Dminus[1807] = 14'b0000000_0000000;
		Dminus[1808] = 14'b0000000_0000000;
		Dminus[1809] = 14'b0000000_0000000;
		Dminus[1810] = 14'b0000000_0000000;
		Dminus[1811] = 14'b0000000_0000000;
		Dminus[1812] = 14'b0000000_0000000;
		Dminus[1813] = 14'b0000000_0000000;
		Dminus[1814] = 14'b0000000_0000000;
		Dminus[1815] = 14'b0000000_0000000;
		Dminus[1816] = 14'b0000000_0000000;
		Dminus[1817] = 14'b0000000_0000000;
		Dminus[1818] = 14'b0000000_0000000;
		Dminus[1819] = 14'b0000000_0000000;
		Dminus[1820] = 14'b0000000_0000000;
		Dminus[1821] = 14'b0000000_0000000;
		Dminus[1822] = 14'b0000000_0000000;
		Dminus[1823] = 14'b0000000_0000000;
		Dminus[1824] = 14'b0000000_0000000;
		Dminus[1825] = 14'b0000000_0000000;
		Dminus[1826] = 14'b0000000_0000000;
		Dminus[1827] = 14'b0000000_0000000;
		Dminus[1828] = 14'b0000000_0000000;
		Dminus[1829] = 14'b0000000_0000000;
		Dminus[1830] = 14'b0000000_0000000;
		Dminus[1831] = 14'b0000000_0000000;
		Dminus[1832] = 14'b0000000_0000000;
		Dminus[1833] = 14'b0000000_0000000;
		Dminus[1834] = 14'b0000000_0000000;
		Dminus[1835] = 14'b0000000_0000000;
		Dminus[1836] = 14'b0000000_0000000;
		Dminus[1837] = 14'b0000000_0000000;
		Dminus[1838] = 14'b0000000_0000000;
		Dminus[1839] = 14'b0000000_0000000;
		Dminus[1840] = 14'b0000000_0000000;
		Dminus[1841] = 14'b0000000_0000000;
		Dminus[1842] = 14'b0000000_0000000;
		Dminus[1843] = 14'b0000000_0000000;
		Dminus[1844] = 14'b0000000_0000000;
		Dminus[1845] = 14'b0000000_0000000;
		Dminus[1846] = 14'b0000000_0000000;
		Dminus[1847] = 14'b0000000_0000000;
		Dminus[1848] = 14'b0000000_0000000;
		Dminus[1849] = 14'b0000000_0000000;
		Dminus[1850] = 14'b0000000_0000000;
		Dminus[1851] = 14'b0000000_0000000;
		Dminus[1852] = 14'b0000000_0000000;
		Dminus[1853] = 14'b0000000_0000000;
		Dminus[1854] = 14'b0000000_0000000;
		Dminus[1855] = 14'b0000000_0000000;
		Dminus[1856] = 14'b0000000_0000000;
		Dminus[1857] = 14'b0000000_0000000;
		Dminus[1858] = 14'b0000000_0000000;
		Dminus[1859] = 14'b0000000_0000000;
		Dminus[1860] = 14'b0000000_0000000;
		Dminus[1861] = 14'b0000000_0000000;
		Dminus[1862] = 14'b0000000_0000000;
		Dminus[1863] = 14'b0000000_0000000;
		Dminus[1864] = 14'b0000000_0000000;
		Dminus[1865] = 14'b0000000_0000000;
		Dminus[1866] = 14'b0000000_0000000;
		Dminus[1867] = 14'b0000000_0000000;
		Dminus[1868] = 14'b0000000_0000000;
		Dminus[1869] = 14'b0000000_0000000;
		Dminus[1870] = 14'b0000000_0000000;
		Dminus[1871] = 14'b0000000_0000000;
		Dminus[1872] = 14'b0000000_0000000;
		Dminus[1873] = 14'b0000000_0000000;
		Dminus[1874] = 14'b0000000_0000000;
		Dminus[1875] = 14'b0000000_0000000;
		Dminus[1876] = 14'b0000000_0000000;
		Dminus[1877] = 14'b0000000_0000000;
		Dminus[1878] = 14'b0000000_0000000;
		Dminus[1879] = 14'b0000000_0000000;
		Dminus[1880] = 14'b0000000_0000000;
		Dminus[1881] = 14'b0000000_0000000;
		Dminus[1882] = 14'b0000000_0000000;
		Dminus[1883] = 14'b0000000_0000000;
		Dminus[1884] = 14'b0000000_0000000;
		Dminus[1885] = 14'b0000000_0000000;
		Dminus[1886] = 14'b0000000_0000000;
		Dminus[1887] = 14'b0000000_0000000;
		Dminus[1888] = 14'b0000000_0000000;
		Dminus[1889] = 14'b0000000_0000000;
		Dminus[1890] = 14'b0000000_0000000;
		Dminus[1891] = 14'b0000000_0000000;
		Dminus[1892] = 14'b0000000_0000000;
		Dminus[1893] = 14'b0000000_0000000;
		Dminus[1894] = 14'b0000000_0000000;
		Dminus[1895] = 14'b0000000_0000000;
		Dminus[1896] = 14'b0000000_0000000;
		Dminus[1897] = 14'b0000000_0000000;
		Dminus[1898] = 14'b0000000_0000000;
		Dminus[1899] = 14'b0000000_0000000;
		Dminus[1900] = 14'b0000000_0000000;
		Dminus[1901] = 14'b0000000_0000000;
		Dminus[1902] = 14'b0000000_0000000;
		Dminus[1903] = 14'b0000000_0000000;
		Dminus[1904] = 14'b0000000_0000000;
		Dminus[1905] = 14'b0000000_0000000;
		Dminus[1906] = 14'b0000000_0000000;
		Dminus[1907] = 14'b0000000_0000000;
		Dminus[1908] = 14'b0000000_0000000;
		Dminus[1909] = 14'b0000000_0000000;
		Dminus[1910] = 14'b0000000_0000000;
		Dminus[1911] = 14'b0000000_0000000;
		Dminus[1912] = 14'b0000000_0000000;
		Dminus[1913] = 14'b0000000_0000000;
		Dminus[1914] = 14'b0000000_0000000;
		Dminus[1915] = 14'b0000000_0000000;
		Dminus[1916] = 14'b0000000_0000000;
		Dminus[1917] = 14'b0000000_0000000;
		Dminus[1918] = 14'b0000000_0000000;
		Dminus[1919] = 14'b0000000_0000000;
		Dminus[1920] = 14'b0000000_0000000;
		Dminus[1921] = 14'b0000000_0000000;
		Dminus[1922] = 14'b0000000_0000000;
		Dminus[1923] = 14'b0000000_0000000;
		Dminus[1924] = 14'b0000000_0000000;
		Dminus[1925] = 14'b0000000_0000000;
		Dminus[1926] = 14'b0000000_0000000;
		Dminus[1927] = 14'b0000000_0000000;
		Dminus[1928] = 14'b0000000_0000000;
		Dminus[1929] = 14'b0000000_0000000;
		Dminus[1930] = 14'b0000000_0000000;
		Dminus[1931] = 14'b0000000_0000000;
		Dminus[1932] = 14'b0000000_0000000;
		Dminus[1933] = 14'b0000000_0000000;
		Dminus[1934] = 14'b0000000_0000000;
		Dminus[1935] = 14'b0000000_0000000;
		Dminus[1936] = 14'b0000000_0000000;
		Dminus[1937] = 14'b0000000_0000000;
		Dminus[1938] = 14'b0000000_0000000;
		Dminus[1939] = 14'b0000000_0000000;
		Dminus[1940] = 14'b0000000_0000000;
		Dminus[1941] = 14'b0000000_0000000;
		Dminus[1942] = 14'b0000000_0000000;
		Dminus[1943] = 14'b0000000_0000000;
		Dminus[1944] = 14'b0000000_0000000;
		Dminus[1945] = 14'b0000000_0000000;
		Dminus[1946] = 14'b0000000_0000000;
		Dminus[1947] = 14'b0000000_0000000;
		Dminus[1948] = 14'b0000000_0000000;
		Dminus[1949] = 14'b0000000_0000000;
		Dminus[1950] = 14'b0000000_0000000;
		Dminus[1951] = 14'b0000000_0000000;
		Dminus[1952] = 14'b0000000_0000000;
		Dminus[1953] = 14'b0000000_0000000;
		Dminus[1954] = 14'b0000000_0000000;
		Dminus[1955] = 14'b0000000_0000000;
		Dminus[1956] = 14'b0000000_0000000;
		Dminus[1957] = 14'b0000000_0000000;
		Dminus[1958] = 14'b0000000_0000000;
		Dminus[1959] = 14'b0000000_0000000;
		Dminus[1960] = 14'b0000000_0000000;
		Dminus[1961] = 14'b0000000_0000000;
		Dminus[1962] = 14'b0000000_0000000;
		Dminus[1963] = 14'b0000000_0000000;
		Dminus[1964] = 14'b0000000_0000000;
		Dminus[1965] = 14'b0000000_0000000;
		Dminus[1966] = 14'b0000000_0000000;
		Dminus[1967] = 14'b0000000_0000000;
		Dminus[1968] = 14'b0000000_0000000;
		Dminus[1969] = 14'b0000000_0000000;
		Dminus[1970] = 14'b0000000_0000000;
		Dminus[1971] = 14'b0000000_0000000;
		Dminus[1972] = 14'b0000000_0000000;
		Dminus[1973] = 14'b0000000_0000000;
		Dminus[1974] = 14'b0000000_0000000;
		Dminus[1975] = 14'b0000000_0000000;
		Dminus[1976] = 14'b0000000_0000000;
		Dminus[1977] = 14'b0000000_0000000;
		Dminus[1978] = 14'b0000000_0000000;
		Dminus[1979] = 14'b0000000_0000000;
		Dminus[1980] = 14'b0000000_0000000;
		Dminus[1981] = 14'b0000000_0000000;
		Dminus[1982] = 14'b0000000_0000000;
		Dminus[1983] = 14'b0000000_0000000;
		Dminus[1984] = 14'b0000000_0000000;
		Dminus[1985] = 14'b0000000_0000000;
		Dminus[1986] = 14'b0000000_0000000;
		Dminus[1987] = 14'b0000000_0000000;
		Dminus[1988] = 14'b0000000_0000000;
		Dminus[1989] = 14'b0000000_0000000;
		Dminus[1990] = 14'b0000000_0000000;
		Dminus[1991] = 14'b0000000_0000000;
		Dminus[1992] = 14'b0000000_0000000;
		Dminus[1993] = 14'b0000000_0000000;
		Dminus[1994] = 14'b0000000_0000000;
		Dminus[1995] = 14'b0000000_0000000;
		Dminus[1996] = 14'b0000000_0000000;
		Dminus[1997] = 14'b0000000_0000000;
		Dminus[1998] = 14'b0000000_0000000;
		Dminus[1999] = 14'b0000000_0000000;
		Dminus[2000] = 14'b0000000_0000000;
		Dminus[2001] = 14'b0000000_0000000;
		Dminus[2002] = 14'b0000000_0000000;
		Dminus[2003] = 14'b0000000_0000000;
		Dminus[2004] = 14'b0000000_0000000;
		Dminus[2005] = 14'b0000000_0000000;
		Dminus[2006] = 14'b0000000_0000000;
		Dminus[2007] = 14'b0000000_0000000;
		Dminus[2008] = 14'b0000000_0000000;
		Dminus[2009] = 14'b0000000_0000000;
		Dminus[2010] = 14'b0000000_0000000;
		Dminus[2011] = 14'b0000000_0000000;
		Dminus[2012] = 14'b0000000_0000000;
		Dminus[2013] = 14'b0000000_0000000;
		Dminus[2014] = 14'b0000000_0000000;
		Dminus[2015] = 14'b0000000_0000000;
		Dminus[2016] = 14'b0000000_0000000;
		Dminus[2017] = 14'b0000000_0000000;
		Dminus[2018] = 14'b0000000_0000000;
		Dminus[2019] = 14'b0000000_0000000;
		Dminus[2020] = 14'b0000000_0000000;
		Dminus[2021] = 14'b0000000_0000000;
		Dminus[2022] = 14'b0000000_0000000;
		Dminus[2023] = 14'b0000000_0000000;
		Dminus[2024] = 14'b0000000_0000000;
		Dminus[2025] = 14'b0000000_0000000;
		Dminus[2026] = 14'b0000000_0000000;
		Dminus[2027] = 14'b0000000_0000000;
		Dminus[2028] = 14'b0000000_0000000;
		Dminus[2029] = 14'b0000000_0000000;
		Dminus[2030] = 14'b0000000_0000000;
		Dminus[2031] = 14'b0000000_0000000;
		Dminus[2032] = 14'b0000000_0000000;
		Dminus[2033] = 14'b0000000_0000000;
		Dminus[2034] = 14'b0000000_0000000;
		Dminus[2035] = 14'b0000000_0000000;
		Dminus[2036] = 14'b0000000_0000000;
		Dminus[2037] = 14'b0000000_0000000;
		Dminus[2038] = 14'b0000000_0000000;
		Dminus[2039] = 14'b0000000_0000000;
		Dminus[2040] = 14'b0000000_0000000;
		Dminus[2041] = 14'b0000000_0000000;
		Dminus[2042] = 14'b0000000_0000000;
		Dminus[2043] = 14'b0000000_0000000;
		Dminus[2044] = 14'b0000000_0000000;
		Dminus[2045] = 14'b0000000_0000000;
		Dminus[2046] = 14'b0000000_0000000;
		Dminus[2047] = 14'b0000000_0000000;
		Dminus[2048] = 14'b0000000_0000000;
		Dminus[2049] = 14'b0000000_0000000;
		Dminus[2050] = 14'b0000000_0000000;
		Dminus[2051] = 14'b0000000_0000000;
		Dminus[2052] = 14'b0000000_0000000;
		Dminus[2053] = 14'b0000000_0000000;
		Dminus[2054] = 14'b0000000_0000000;
		Dminus[2055] = 14'b0000000_0000000;
		Dminus[2056] = 14'b0000000_0000000;
		Dminus[2057] = 14'b0000000_0000000;
		Dminus[2058] = 14'b0000000_0000000;
		Dminus[2059] = 14'b0000000_0000000;
		Dminus[2060] = 14'b0000000_0000000;
		Dminus[2061] = 14'b0000000_0000000;
		Dminus[2062] = 14'b0000000_0000000;
		Dminus[2063] = 14'b0000000_0000000;
		Dminus[2064] = 14'b0000000_0000000;
		Dminus[2065] = 14'b0000000_0000000;
		Dminus[2066] = 14'b0000000_0000000;
		Dminus[2067] = 14'b0000000_0000000;
		Dminus[2068] = 14'b0000000_0000000;
		Dminus[2069] = 14'b0000000_0000000;
		Dminus[2070] = 14'b0000000_0000000;
		Dminus[2071] = 14'b0000000_0000000;
		Dminus[2072] = 14'b0000000_0000000;
		Dminus[2073] = 14'b0000000_0000000;
		Dminus[2074] = 14'b0000000_0000000;
		Dminus[2075] = 14'b0000000_0000000;
		Dminus[2076] = 14'b0000000_0000000;
		Dminus[2077] = 14'b0000000_0000000;
		Dminus[2078] = 14'b0000000_0000000;
		Dminus[2079] = 14'b0000000_0000000;
		Dminus[2080] = 14'b0000000_0000000;
		Dminus[2081] = 14'b0000000_0000000;
		Dminus[2082] = 14'b0000000_0000000;
		Dminus[2083] = 14'b0000000_0000000;
		Dminus[2084] = 14'b0000000_0000000;
		Dminus[2085] = 14'b0000000_0000000;
		Dminus[2086] = 14'b0000000_0000000;
		Dminus[2087] = 14'b0000000_0000000;
		Dminus[2088] = 14'b0000000_0000000;
		Dminus[2089] = 14'b0000000_0000000;
		Dminus[2090] = 14'b0000000_0000000;
		Dminus[2091] = 14'b0000000_0000000;
		Dminus[2092] = 14'b0000000_0000000;
		Dminus[2093] = 14'b0000000_0000000;
		Dminus[2094] = 14'b0000000_0000000;
		Dminus[2095] = 14'b0000000_0000000;
		Dminus[2096] = 14'b0000000_0000000;
		Dminus[2097] = 14'b0000000_0000000;
		Dminus[2098] = 14'b0000000_0000000;
		Dminus[2099] = 14'b0000000_0000000;
		Dminus[2100] = 14'b0000000_0000000;
		Dminus[2101] = 14'b0000000_0000000;
		Dminus[2102] = 14'b0000000_0000000;
		Dminus[2103] = 14'b0000000_0000000;
		Dminus[2104] = 14'b0000000_0000000;
		Dminus[2105] = 14'b0000000_0000000;
		Dminus[2106] = 14'b0000000_0000000;
		Dminus[2107] = 14'b0000000_0000000;
		Dminus[2108] = 14'b0000000_0000000;
		Dminus[2109] = 14'b0000000_0000000;
		Dminus[2110] = 14'b0000000_0000000;
		Dminus[2111] = 14'b0000000_0000000;
		Dminus[2112] = 14'b0000000_0000000;
		Dminus[2113] = 14'b0000000_0000000;
		Dminus[2114] = 14'b0000000_0000000;
		Dminus[2115] = 14'b0000000_0000000;
		Dminus[2116] = 14'b0000000_0000000;
		Dminus[2117] = 14'b0000000_0000000;
		Dminus[2118] = 14'b0000000_0000000;
		Dminus[2119] = 14'b0000000_0000000;
		Dminus[2120] = 14'b0000000_0000000;
		Dminus[2121] = 14'b0000000_0000000;
		Dminus[2122] = 14'b0000000_0000000;
		Dminus[2123] = 14'b0000000_0000000;
		Dminus[2124] = 14'b0000000_0000000;
		Dminus[2125] = 14'b0000000_0000000;
		Dminus[2126] = 14'b0000000_0000000;
		Dminus[2127] = 14'b0000000_0000000;
		Dminus[2128] = 14'b0000000_0000000;
		Dminus[2129] = 14'b0000000_0000000;
		Dminus[2130] = 14'b0000000_0000000;
		Dminus[2131] = 14'b0000000_0000000;
		Dminus[2132] = 14'b0000000_0000000;
		Dminus[2133] = 14'b0000000_0000000;
		Dminus[2134] = 14'b0000000_0000000;
		Dminus[2135] = 14'b0000000_0000000;
		Dminus[2136] = 14'b0000000_0000000;
		Dminus[2137] = 14'b0000000_0000000;
		Dminus[2138] = 14'b0000000_0000000;
		Dminus[2139] = 14'b0000000_0000000;
		Dminus[2140] = 14'b0000000_0000000;
		Dminus[2141] = 14'b0000000_0000000;
		Dminus[2142] = 14'b0000000_0000000;
		Dminus[2143] = 14'b0000000_0000000;
		Dminus[2144] = 14'b0000000_0000000;
		Dminus[2145] = 14'b0000000_0000000;
		Dminus[2146] = 14'b0000000_0000000;
		Dminus[2147] = 14'b0000000_0000000;
		Dminus[2148] = 14'b0000000_0000000;
		Dminus[2149] = 14'b0000000_0000000;
		Dminus[2150] = 14'b0000000_0000000;
		Dminus[2151] = 14'b0000000_0000000;
		Dminus[2152] = 14'b0000000_0000000;
		Dminus[2153] = 14'b0000000_0000000;
		Dminus[2154] = 14'b0000000_0000000;
		Dminus[2155] = 14'b0000000_0000000;
		Dminus[2156] = 14'b0000000_0000000;
		Dminus[2157] = 14'b0000000_0000000;
		Dminus[2158] = 14'b0000000_0000000;
		Dminus[2159] = 14'b0000000_0000000;
		Dminus[2160] = 14'b0000000_0000000;
		Dminus[2161] = 14'b0000000_0000000;
		Dminus[2162] = 14'b0000000_0000000;
		Dminus[2163] = 14'b0000000_0000000;
		Dminus[2164] = 14'b0000000_0000000;
		Dminus[2165] = 14'b0000000_0000000;
		Dminus[2166] = 14'b0000000_0000000;
		Dminus[2167] = 14'b0000000_0000000;
		Dminus[2168] = 14'b0000000_0000000;
		Dminus[2169] = 14'b0000000_0000000;
		Dminus[2170] = 14'b0000000_0000000;
		Dminus[2171] = 14'b0000000_0000000;
		Dminus[2172] = 14'b0000000_0000000;
		Dminus[2173] = 14'b0000000_0000000;
		Dminus[2174] = 14'b0000000_0000000;
		Dminus[2175] = 14'b0000000_0000000;
		Dminus[2176] = 14'b0000000_0000000;
		Dminus[2177] = 14'b0000000_0000000;
		Dminus[2178] = 14'b0000000_0000000;
		Dminus[2179] = 14'b0000000_0000000;
		Dminus[2180] = 14'b0000000_0000000;
		Dminus[2181] = 14'b0000000_0000000;
		Dminus[2182] = 14'b0000000_0000000;
		Dminus[2183] = 14'b0000000_0000000;
		Dminus[2184] = 14'b0000000_0000000;
		Dminus[2185] = 14'b0000000_0000000;
		Dminus[2186] = 14'b0000000_0000000;
		Dminus[2187] = 14'b0000000_0000000;
		Dminus[2188] = 14'b0000000_0000000;
		Dminus[2189] = 14'b0000000_0000000;
		Dminus[2190] = 14'b0000000_0000000;
		Dminus[2191] = 14'b0000000_0000000;
		Dminus[2192] = 14'b0000000_0000000;
		Dminus[2193] = 14'b0000000_0000000;
		Dminus[2194] = 14'b0000000_0000000;
		Dminus[2195] = 14'b0000000_0000000;
		Dminus[2196] = 14'b0000000_0000000;
		Dminus[2197] = 14'b0000000_0000000;
		Dminus[2198] = 14'b0000000_0000000;
		Dminus[2199] = 14'b0000000_0000000;
		Dminus[2200] = 14'b0000000_0000000;
		Dminus[2201] = 14'b0000000_0000000;
		Dminus[2202] = 14'b0000000_0000000;
		Dminus[2203] = 14'b0000000_0000000;
		Dminus[2204] = 14'b0000000_0000000;
		Dminus[2205] = 14'b0000000_0000000;
		Dminus[2206] = 14'b0000000_0000000;
		Dminus[2207] = 14'b0000000_0000000;
		Dminus[2208] = 14'b0000000_0000000;
		Dminus[2209] = 14'b0000000_0000000;
		Dminus[2210] = 14'b0000000_0000000;
		Dminus[2211] = 14'b0000000_0000000;
		Dminus[2212] = 14'b0000000_0000000;
		Dminus[2213] = 14'b0000000_0000000;
		Dminus[2214] = 14'b0000000_0000000;
		Dminus[2215] = 14'b0000000_0000000;
		Dminus[2216] = 14'b0000000_0000000;
		Dminus[2217] = 14'b0000000_0000000;
		Dminus[2218] = 14'b0000000_0000000;
		Dminus[2219] = 14'b0000000_0000000;
		Dminus[2220] = 14'b0000000_0000000;
		Dminus[2221] = 14'b0000000_0000000;
		Dminus[2222] = 14'b0000000_0000000;
		Dminus[2223] = 14'b0000000_0000000;
		Dminus[2224] = 14'b0000000_0000000;
		Dminus[2225] = 14'b0000000_0000000;
		Dminus[2226] = 14'b0000000_0000000;
		Dminus[2227] = 14'b0000000_0000000;
		Dminus[2228] = 14'b0000000_0000000;
		Dminus[2229] = 14'b0000000_0000000;
		Dminus[2230] = 14'b0000000_0000000;
		Dminus[2231] = 14'b0000000_0000000;
		Dminus[2232] = 14'b0000000_0000000;
		Dminus[2233] = 14'b0000000_0000000;
		Dminus[2234] = 14'b0000000_0000000;
		Dminus[2235] = 14'b0000000_0000000;
		Dminus[2236] = 14'b0000000_0000000;
		Dminus[2237] = 14'b0000000_0000000;
		Dminus[2238] = 14'b0000000_0000000;
		Dminus[2239] = 14'b0000000_0000000;
		Dminus[2240] = 14'b0000000_0000000;
		Dminus[2241] = 14'b0000000_0000000;
		Dminus[2242] = 14'b0000000_0000000;
		Dminus[2243] = 14'b0000000_0000000;
		Dminus[2244] = 14'b0000000_0000000;
		Dminus[2245] = 14'b0000000_0000000;
		Dminus[2246] = 14'b0000000_0000000;
		Dminus[2247] = 14'b0000000_0000000;
		Dminus[2248] = 14'b0000000_0000000;
		Dminus[2249] = 14'b0000000_0000000;
		Dminus[2250] = 14'b0000000_0000000;
		Dminus[2251] = 14'b0000000_0000000;
		Dminus[2252] = 14'b0000000_0000000;
		Dminus[2253] = 14'b0000000_0000000;
		Dminus[2254] = 14'b0000000_0000000;
		Dminus[2255] = 14'b0000000_0000000;
		Dminus[2256] = 14'b0000000_0000000;
		Dminus[2257] = 14'b0000000_0000000;
		Dminus[2258] = 14'b0000000_0000000;
		Dminus[2259] = 14'b0000000_0000000;
		Dminus[2260] = 14'b0000000_0000000;
		Dminus[2261] = 14'b0000000_0000000;
		Dminus[2262] = 14'b0000000_0000000;
		Dminus[2263] = 14'b0000000_0000000;
		Dminus[2264] = 14'b0000000_0000000;
		Dminus[2265] = 14'b0000000_0000000;
		Dminus[2266] = 14'b0000000_0000000;
		Dminus[2267] = 14'b0000000_0000000;
		Dminus[2268] = 14'b0000000_0000000;
		Dminus[2269] = 14'b0000000_0000000;
		Dminus[2270] = 14'b0000000_0000000;
		Dminus[2271] = 14'b0000000_0000000;
		Dminus[2272] = 14'b0000000_0000000;
		Dminus[2273] = 14'b0000000_0000000;
		Dminus[2274] = 14'b0000000_0000000;
		Dminus[2275] = 14'b0000000_0000000;
		Dminus[2276] = 14'b0000000_0000000;
		Dminus[2277] = 14'b0000000_0000000;
		Dminus[2278] = 14'b0000000_0000000;
		Dminus[2279] = 14'b0000000_0000000;
		Dminus[2280] = 14'b0000000_0000000;
		Dminus[2281] = 14'b0000000_0000000;
		Dminus[2282] = 14'b0000000_0000000;
		Dminus[2283] = 14'b0000000_0000000;
		Dminus[2284] = 14'b0000000_0000000;
		Dminus[2285] = 14'b0000000_0000000;
		Dminus[2286] = 14'b0000000_0000000;
		Dminus[2287] = 14'b0000000_0000000;
		Dminus[2288] = 14'b0000000_0000000;
		Dminus[2289] = 14'b0000000_0000000;
		Dminus[2290] = 14'b0000000_0000000;
		Dminus[2291] = 14'b0000000_0000000;
		Dminus[2292] = 14'b0000000_0000000;
		Dminus[2293] = 14'b0000000_0000000;
		Dminus[2294] = 14'b0000000_0000000;
		Dminus[2295] = 14'b0000000_0000000;
		Dminus[2296] = 14'b0000000_0000000;
		Dminus[2297] = 14'b0000000_0000000;
		Dminus[2298] = 14'b0000000_0000000;
		Dminus[2299] = 14'b0000000_0000000;
		Dminus[2300] = 14'b0000000_0000000;
		Dminus[2301] = 14'b0000000_0000000;
		Dminus[2302] = 14'b0000000_0000000;
		Dminus[2303] = 14'b0000000_0000000;
		Dminus[2304] = 14'b0000000_0000000;
		Dminus[2305] = 14'b0000000_0000000;
		Dminus[2306] = 14'b0000000_0000000;
		Dminus[2307] = 14'b0000000_0000000;
		Dminus[2308] = 14'b0000000_0000000;
		Dminus[2309] = 14'b0000000_0000000;
		Dminus[2310] = 14'b0000000_0000000;
		Dminus[2311] = 14'b0000000_0000000;
		Dminus[2312] = 14'b0000000_0000000;
		Dminus[2313] = 14'b0000000_0000000;
		Dminus[2314] = 14'b0000000_0000000;
		Dminus[2315] = 14'b0000000_0000000;
		Dminus[2316] = 14'b0000000_0000000;
		Dminus[2317] = 14'b0000000_0000000;
		Dminus[2318] = 14'b0000000_0000000;
		Dminus[2319] = 14'b0000000_0000000;
		Dminus[2320] = 14'b0000000_0000000;
		Dminus[2321] = 14'b0000000_0000000;
		Dminus[2322] = 14'b0000000_0000000;
		Dminus[2323] = 14'b0000000_0000000;
		Dminus[2324] = 14'b0000000_0000000;
		Dminus[2325] = 14'b0000000_0000000;
		Dminus[2326] = 14'b0000000_0000000;
		Dminus[2327] = 14'b0000000_0000000;
		Dminus[2328] = 14'b0000000_0000000;
		Dminus[2329] = 14'b0000000_0000000;
		Dminus[2330] = 14'b0000000_0000000;
		Dminus[2331] = 14'b0000000_0000000;
		Dminus[2332] = 14'b0000000_0000000;
		Dminus[2333] = 14'b0000000_0000000;
		Dminus[2334] = 14'b0000000_0000000;
		Dminus[2335] = 14'b0000000_0000000;
		Dminus[2336] = 14'b0000000_0000000;
		Dminus[2337] = 14'b0000000_0000000;
		Dminus[2338] = 14'b0000000_0000000;
		Dminus[2339] = 14'b0000000_0000000;
		Dminus[2340] = 14'b0000000_0000000;
		Dminus[2341] = 14'b0000000_0000000;
		Dminus[2342] = 14'b0000000_0000000;
		Dminus[2343] = 14'b0000000_0000000;
		Dminus[2344] = 14'b0000000_0000000;
		Dminus[2345] = 14'b0000000_0000000;
		Dminus[2346] = 14'b0000000_0000000;
		Dminus[2347] = 14'b0000000_0000000;
		Dminus[2348] = 14'b0000000_0000000;
		Dminus[2349] = 14'b0000000_0000000;
		Dminus[2350] = 14'b0000000_0000000;
		Dminus[2351] = 14'b0000000_0000000;
		Dminus[2352] = 14'b0000000_0000000;
		Dminus[2353] = 14'b0000000_0000000;
		Dminus[2354] = 14'b0000000_0000000;
		Dminus[2355] = 14'b0000000_0000000;
		Dminus[2356] = 14'b0000000_0000000;
		Dminus[2357] = 14'b0000000_0000000;
		Dminus[2358] = 14'b0000000_0000000;
		Dminus[2359] = 14'b0000000_0000000;
		Dminus[2360] = 14'b0000000_0000000;
		Dminus[2361] = 14'b0000000_0000000;
		Dminus[2362] = 14'b0000000_0000000;
		Dminus[2363] = 14'b0000000_0000000;
		Dminus[2364] = 14'b0000000_0000000;
		Dminus[2365] = 14'b0000000_0000000;
		Dminus[2366] = 14'b0000000_0000000;
		Dminus[2367] = 14'b0000000_0000000;
		Dminus[2368] = 14'b0000000_0000000;
		Dminus[2369] = 14'b0000000_0000000;
		Dminus[2370] = 14'b0000000_0000000;
		Dminus[2371] = 14'b0000000_0000000;
		Dminus[2372] = 14'b0000000_0000000;
		Dminus[2373] = 14'b0000000_0000000;
		Dminus[2374] = 14'b0000000_0000000;
		Dminus[2375] = 14'b0000000_0000000;
		Dminus[2376] = 14'b0000000_0000000;
		Dminus[2377] = 14'b0000000_0000000;
		Dminus[2378] = 14'b0000000_0000000;
		Dminus[2379] = 14'b0000000_0000000;
		Dminus[2380] = 14'b0000000_0000000;
		Dminus[2381] = 14'b0000000_0000000;
		Dminus[2382] = 14'b0000000_0000000;
		Dminus[2383] = 14'b0000000_0000000;
		Dminus[2384] = 14'b0000000_0000000;
		Dminus[2385] = 14'b0000000_0000000;
		Dminus[2386] = 14'b0000000_0000000;
		Dminus[2387] = 14'b0000000_0000000;
		Dminus[2388] = 14'b0000000_0000000;
		Dminus[2389] = 14'b0000000_0000000;
		Dminus[2390] = 14'b0000000_0000000;
		Dminus[2391] = 14'b0000000_0000000;
		Dminus[2392] = 14'b0000000_0000000;
		Dminus[2393] = 14'b0000000_0000000;
		Dminus[2394] = 14'b0000000_0000000;
		Dminus[2395] = 14'b0000000_0000000;
		Dminus[2396] = 14'b0000000_0000000;
		Dminus[2397] = 14'b0000000_0000000;
		Dminus[2398] = 14'b0000000_0000000;
		Dminus[2399] = 14'b0000000_0000000;
		Dminus[2400] = 14'b0000000_0000000;
		Dminus[2401] = 14'b0000000_0000000;
		Dminus[2402] = 14'b0000000_0000000;
		Dminus[2403] = 14'b0000000_0000000;
		Dminus[2404] = 14'b0000000_0000000;
		Dminus[2405] = 14'b0000000_0000000;
		Dminus[2406] = 14'b0000000_0000000;
		Dminus[2407] = 14'b0000000_0000000;
		Dminus[2408] = 14'b0000000_0000000;
		Dminus[2409] = 14'b0000000_0000000;
		Dminus[2410] = 14'b0000000_0000000;
		Dminus[2411] = 14'b0000000_0000000;
		Dminus[2412] = 14'b0000000_0000000;
		Dminus[2413] = 14'b0000000_0000000;
		Dminus[2414] = 14'b0000000_0000000;
		Dminus[2415] = 14'b0000000_0000000;
		Dminus[2416] = 14'b0000000_0000000;
		Dminus[2417] = 14'b0000000_0000000;
		Dminus[2418] = 14'b0000000_0000000;
		Dminus[2419] = 14'b0000000_0000000;
		Dminus[2420] = 14'b0000000_0000000;
		Dminus[2421] = 14'b0000000_0000000;
		Dminus[2422] = 14'b0000000_0000000;
		Dminus[2423] = 14'b0000000_0000000;
		Dminus[2424] = 14'b0000000_0000000;
		Dminus[2425] = 14'b0000000_0000000;
		Dminus[2426] = 14'b0000000_0000000;
		Dminus[2427] = 14'b0000000_0000000;
		Dminus[2428] = 14'b0000000_0000000;
		Dminus[2429] = 14'b0000000_0000000;
		Dminus[2430] = 14'b0000000_0000000;
		Dminus[2431] = 14'b0000000_0000000;
		Dminus[2432] = 14'b0000000_0000000;
		Dminus[2433] = 14'b0000000_0000000;
		Dminus[2434] = 14'b0000000_0000000;
		Dminus[2435] = 14'b0000000_0000000;
		Dminus[2436] = 14'b0000000_0000000;
		Dminus[2437] = 14'b0000000_0000000;
		Dminus[2438] = 14'b0000000_0000000;
		Dminus[2439] = 14'b0000000_0000000;
		Dminus[2440] = 14'b0000000_0000000;
		Dminus[2441] = 14'b0000000_0000000;
		Dminus[2442] = 14'b0000000_0000000;
		Dminus[2443] = 14'b0000000_0000000;
		Dminus[2444] = 14'b0000000_0000000;
		Dminus[2445] = 14'b0000000_0000000;
		Dminus[2446] = 14'b0000000_0000000;
		Dminus[2447] = 14'b0000000_0000000;
		Dminus[2448] = 14'b0000000_0000000;
		Dminus[2449] = 14'b0000000_0000000;
		Dminus[2450] = 14'b0000000_0000000;
		Dminus[2451] = 14'b0000000_0000000;
		Dminus[2452] = 14'b0000000_0000000;
		Dminus[2453] = 14'b0000000_0000000;
		Dminus[2454] = 14'b0000000_0000000;
		Dminus[2455] = 14'b0000000_0000000;
		Dminus[2456] = 14'b0000000_0000000;
		Dminus[2457] = 14'b0000000_0000000;
		Dminus[2458] = 14'b0000000_0000000;
		Dminus[2459] = 14'b0000000_0000000;
		Dminus[2460] = 14'b0000000_0000000;
		Dminus[2461] = 14'b0000000_0000000;
		Dminus[2462] = 14'b0000000_0000000;
		Dminus[2463] = 14'b0000000_0000000;
		Dminus[2464] = 14'b0000000_0000000;
		Dminus[2465] = 14'b0000000_0000000;
		Dminus[2466] = 14'b0000000_0000000;
		Dminus[2467] = 14'b0000000_0000000;
		Dminus[2468] = 14'b0000000_0000000;
		Dminus[2469] = 14'b0000000_0000000;
		Dminus[2470] = 14'b0000000_0000000;
		Dminus[2471] = 14'b0000000_0000000;
		Dminus[2472] = 14'b0000000_0000000;
		Dminus[2473] = 14'b0000000_0000000;
		Dminus[2474] = 14'b0000000_0000000;
		Dminus[2475] = 14'b0000000_0000000;
		Dminus[2476] = 14'b0000000_0000000;
		Dminus[2477] = 14'b0000000_0000000;
		Dminus[2478] = 14'b0000000_0000000;
		Dminus[2479] = 14'b0000000_0000000;
		Dminus[2480] = 14'b0000000_0000000;
		Dminus[2481] = 14'b0000000_0000000;
		Dminus[2482] = 14'b0000000_0000000;
		Dminus[2483] = 14'b0000000_0000000;
		Dminus[2484] = 14'b0000000_0000000;
		Dminus[2485] = 14'b0000000_0000000;
		Dminus[2486] = 14'b0000000_0000000;
		Dminus[2487] = 14'b0000000_0000000;
		Dminus[2488] = 14'b0000000_0000000;
		Dminus[2489] = 14'b0000000_0000000;
		Dminus[2490] = 14'b0000000_0000000;
		Dminus[2491] = 14'b0000000_0000000;
		Dminus[2492] = 14'b0000000_0000000;
		Dminus[2493] = 14'b0000000_0000000;
		Dminus[2494] = 14'b0000000_0000000;
		Dminus[2495] = 14'b0000000_0000000;
		Dminus[2496] = 14'b0000000_0000000;
		Dminus[2497] = 14'b0000000_0000000;
		Dminus[2498] = 14'b0000000_0000000;
		Dminus[2499] = 14'b0000000_0000000;
		Dminus[2500] = 14'b0000000_0000000;
		Dminus[2501] = 14'b0000000_0000000;
		Dminus[2502] = 14'b0000000_0000000;
		Dminus[2503] = 14'b0000000_0000000;
		Dminus[2504] = 14'b0000000_0000000;
		Dminus[2505] = 14'b0000000_0000000;
		Dminus[2506] = 14'b0000000_0000000;
		Dminus[2507] = 14'b0000000_0000000;
		Dminus[2508] = 14'b0000000_0000000;
		Dminus[2509] = 14'b0000000_0000000;
		Dminus[2510] = 14'b0000000_0000000;
		Dminus[2511] = 14'b0000000_0000000;
		Dminus[2512] = 14'b0000000_0000000;
		Dminus[2513] = 14'b0000000_0000000;
		Dminus[2514] = 14'b0000000_0000000;
		Dminus[2515] = 14'b0000000_0000000;
		Dminus[2516] = 14'b0000000_0000000;
		Dminus[2517] = 14'b0000000_0000000;
		Dminus[2518] = 14'b0000000_0000000;
		Dminus[2519] = 14'b0000000_0000000;
		Dminus[2520] = 14'b0000000_0000000;
		Dminus[2521] = 14'b0000000_0000000;
		Dminus[2522] = 14'b0000000_0000000;
		Dminus[2523] = 14'b0000000_0000000;
		Dminus[2524] = 14'b0000000_0000000;
		Dminus[2525] = 14'b0000000_0000000;
		Dminus[2526] = 14'b0000000_0000000;
		Dminus[2527] = 14'b0000000_0000000;
		Dminus[2528] = 14'b0000000_0000000;
		Dminus[2529] = 14'b0000000_0000000;
		Dminus[2530] = 14'b0000000_0000000;
		Dminus[2531] = 14'b0000000_0000000;
		Dminus[2532] = 14'b0000000_0000000;
		Dminus[2533] = 14'b0000000_0000000;
		Dminus[2534] = 14'b0000000_0000000;
		Dminus[2535] = 14'b0000000_0000000;
		Dminus[2536] = 14'b0000000_0000000;
		Dminus[2537] = 14'b0000000_0000000;
		Dminus[2538] = 14'b0000000_0000000;
		Dminus[2539] = 14'b0000000_0000000;
		Dminus[2540] = 14'b0000000_0000000;
		Dminus[2541] = 14'b0000000_0000000;
		Dminus[2542] = 14'b0000000_0000000;
		Dminus[2543] = 14'b0000000_0000000;
		Dminus[2544] = 14'b0000000_0000000;
		Dminus[2545] = 14'b0000000_0000000;
		Dminus[2546] = 14'b0000000_0000000;
		Dminus[2547] = 14'b0000000_0000000;
		Dminus[2548] = 14'b0000000_0000000;
		Dminus[2549] = 14'b0000000_0000000;
		Dminus[2550] = 14'b0000000_0000000;
		Dminus[2551] = 14'b0000000_0000000;
		Dminus[2552] = 14'b0000000_0000000;
		Dminus[2553] = 14'b0000000_0000000;
		Dminus[2554] = 14'b0000000_0000000;
		Dminus[2555] = 14'b0000000_0000000;
		Dminus[2556] = 14'b0000000_0000000;
		Dminus[2557] = 14'b0000000_0000000;
		Dminus[2558] = 14'b0000000_0000000;
		Dminus[2559] = 14'b0000000_0000000;
		Dminus[2560] = 14'b0000000_0000000;
		Dminus[2561] = 14'b0000000_0000000;
		Dminus[2562] = 14'b0000000_0000000;
		Dminus[2563] = 14'b0000000_0000000;
		Dminus[2564] = 14'b0000000_0000000;
		Dminus[2565] = 14'b0000000_0000000;
		Dminus[2566] = 14'b0000000_0000000;
		Dminus[2567] = 14'b0000000_0000000;
		Dminus[2568] = 14'b0000000_0000000;
		Dminus[2569] = 14'b0000000_0000000;
		Dminus[2570] = 14'b0000000_0000000;
		Dminus[2571] = 14'b0000000_0000000;
		Dminus[2572] = 14'b0000000_0000000;
		Dminus[2573] = 14'b0000000_0000000;
		Dminus[2574] = 14'b0000000_0000000;
		Dminus[2575] = 14'b0000000_0000000;
		Dminus[2576] = 14'b0000000_0000000;
		Dminus[2577] = 14'b0000000_0000000;
		Dminus[2578] = 14'b0000000_0000000;
		Dminus[2579] = 14'b0000000_0000000;
		Dminus[2580] = 14'b0000000_0000000;
		Dminus[2581] = 14'b0000000_0000000;
		Dminus[2582] = 14'b0000000_0000000;
		Dminus[2583] = 14'b0000000_0000000;
		Dminus[2584] = 14'b0000000_0000000;
		Dminus[2585] = 14'b0000000_0000000;
		Dminus[2586] = 14'b0000000_0000000;
		Dminus[2587] = 14'b0000000_0000000;
		Dminus[2588] = 14'b0000000_0000000;
		Dminus[2589] = 14'b0000000_0000000;
		Dminus[2590] = 14'b0000000_0000000;
		Dminus[2591] = 14'b0000000_0000000;
		Dminus[2592] = 14'b0000000_0000000;
		Dminus[2593] = 14'b0000000_0000000;
		Dminus[2594] = 14'b0000000_0000000;
		Dminus[2595] = 14'b0000000_0000000;
		Dminus[2596] = 14'b0000000_0000000;
		Dminus[2597] = 14'b0000000_0000000;
		Dminus[2598] = 14'b0000000_0000000;
		Dminus[2599] = 14'b0000000_0000000;
		Dminus[2600] = 14'b0000000_0000000;
		Dminus[2601] = 14'b0000000_0000000;
		Dminus[2602] = 14'b0000000_0000000;
		Dminus[2603] = 14'b0000000_0000000;
		Dminus[2604] = 14'b0000000_0000000;
		Dminus[2605] = 14'b0000000_0000000;
		Dminus[2606] = 14'b0000000_0000000;
		Dminus[2607] = 14'b0000000_0000000;
		Dminus[2608] = 14'b0000000_0000000;
		Dminus[2609] = 14'b0000000_0000000;
		Dminus[2610] = 14'b0000000_0000000;
		Dminus[2611] = 14'b0000000_0000000;
		Dminus[2612] = 14'b0000000_0000000;
		Dminus[2613] = 14'b0000000_0000000;
		Dminus[2614] = 14'b0000000_0000000;
		Dminus[2615] = 14'b0000000_0000000;
		Dminus[2616] = 14'b0000000_0000000;
		Dminus[2617] = 14'b0000000_0000000;
		Dminus[2618] = 14'b0000000_0000000;
		Dminus[2619] = 14'b0000000_0000000;
		Dminus[2620] = 14'b0000000_0000000;
		Dminus[2621] = 14'b0000000_0000000;
		Dminus[2622] = 14'b0000000_0000000;
		Dminus[2623] = 14'b0000000_0000000;
		Dminus[2624] = 14'b0000000_0000000;
		Dminus[2625] = 14'b0000000_0000000;
		Dminus[2626] = 14'b0000000_0000000;
		Dminus[2627] = 14'b0000000_0000000;
		Dminus[2628] = 14'b0000000_0000000;
		Dminus[2629] = 14'b0000000_0000000;
		Dminus[2630] = 14'b0000000_0000000;
		Dminus[2631] = 14'b0000000_0000000;
		Dminus[2632] = 14'b0000000_0000000;
		Dminus[2633] = 14'b0000000_0000000;
		Dminus[2634] = 14'b0000000_0000000;
		Dminus[2635] = 14'b0000000_0000000;
		Dminus[2636] = 14'b0000000_0000000;
		Dminus[2637] = 14'b0000000_0000000;
		Dminus[2638] = 14'b0000000_0000000;
		Dminus[2639] = 14'b0000000_0000000;
		Dminus[2640] = 14'b0000000_0000000;
		Dminus[2641] = 14'b0000000_0000000;
		Dminus[2642] = 14'b0000000_0000000;
		Dminus[2643] = 14'b0000000_0000000;
		Dminus[2644] = 14'b0000000_0000000;
		Dminus[2645] = 14'b0000000_0000000;
		Dminus[2646] = 14'b0000000_0000000;
		Dminus[2647] = 14'b0000000_0000000;
		Dminus[2648] = 14'b0000000_0000000;
		Dminus[2649] = 14'b0000000_0000000;
		Dminus[2650] = 14'b0000000_0000000;
		Dminus[2651] = 14'b0000000_0000000;
		Dminus[2652] = 14'b0000000_0000000;
		Dminus[2653] = 14'b0000000_0000000;
		Dminus[2654] = 14'b0000000_0000000;
		Dminus[2655] = 14'b0000000_0000000;
		Dminus[2656] = 14'b0000000_0000000;
		Dminus[2657] = 14'b0000000_0000000;
		Dminus[2658] = 14'b0000000_0000000;
		Dminus[2659] = 14'b0000000_0000000;
		Dminus[2660] = 14'b0000000_0000000;
		Dminus[2661] = 14'b0000000_0000000;
		Dminus[2662] = 14'b0000000_0000000;
		Dminus[2663] = 14'b0000000_0000000;
		Dminus[2664] = 14'b0000000_0000000;
		Dminus[2665] = 14'b0000000_0000000;
		Dminus[2666] = 14'b0000000_0000000;
		Dminus[2667] = 14'b0000000_0000000;
		Dminus[2668] = 14'b0000000_0000000;
		Dminus[2669] = 14'b0000000_0000000;
		Dminus[2670] = 14'b0000000_0000000;
		Dminus[2671] = 14'b0000000_0000000;
		Dminus[2672] = 14'b0000000_0000000;
		Dminus[2673] = 14'b0000000_0000000;
		Dminus[2674] = 14'b0000000_0000000;
		Dminus[2675] = 14'b0000000_0000000;
		Dminus[2676] = 14'b0000000_0000000;
		Dminus[2677] = 14'b0000000_0000000;
		Dminus[2678] = 14'b0000000_0000000;
		Dminus[2679] = 14'b0000000_0000000;
		Dminus[2680] = 14'b0000000_0000000;
		Dminus[2681] = 14'b0000000_0000000;
		Dminus[2682] = 14'b0000000_0000000;
		Dminus[2683] = 14'b0000000_0000000;
		Dminus[2684] = 14'b0000000_0000000;
		Dminus[2685] = 14'b0000000_0000000;
		Dminus[2686] = 14'b0000000_0000000;
		Dminus[2687] = 14'b0000000_0000000;
		Dminus[2688] = 14'b0000000_0000000;
		Dminus[2689] = 14'b0000000_0000000;
		Dminus[2690] = 14'b0000000_0000000;
		Dminus[2691] = 14'b0000000_0000000;
		Dminus[2692] = 14'b0000000_0000000;
		Dminus[2693] = 14'b0000000_0000000;
		Dminus[2694] = 14'b0000000_0000000;
		Dminus[2695] = 14'b0000000_0000000;
		Dminus[2696] = 14'b0000000_0000000;
		Dminus[2697] = 14'b0000000_0000000;
		Dminus[2698] = 14'b0000000_0000000;
		Dminus[2699] = 14'b0000000_0000000;
		Dminus[2700] = 14'b0000000_0000000;
		Dminus[2701] = 14'b0000000_0000000;
		Dminus[2702] = 14'b0000000_0000000;
		Dminus[2703] = 14'b0000000_0000000;
		Dminus[2704] = 14'b0000000_0000000;
		Dminus[2705] = 14'b0000000_0000000;
		Dminus[2706] = 14'b0000000_0000000;
		Dminus[2707] = 14'b0000000_0000000;
		Dminus[2708] = 14'b0000000_0000000;
		Dminus[2709] = 14'b0000000_0000000;
		Dminus[2710] = 14'b0000000_0000000;
		Dminus[2711] = 14'b0000000_0000000;
		Dminus[2712] = 14'b0000000_0000000;
		Dminus[2713] = 14'b0000000_0000000;
		Dminus[2714] = 14'b0000000_0000000;
		Dminus[2715] = 14'b0000000_0000000;
		Dminus[2716] = 14'b0000000_0000000;
		Dminus[2717] = 14'b0000000_0000000;
		Dminus[2718] = 14'b0000000_0000000;
		Dminus[2719] = 14'b0000000_0000000;
		Dminus[2720] = 14'b0000000_0000000;
		Dminus[2721] = 14'b0000000_0000000;
		Dminus[2722] = 14'b0000000_0000000;
		Dminus[2723] = 14'b0000000_0000000;
		Dminus[2724] = 14'b0000000_0000000;
		Dminus[2725] = 14'b0000000_0000000;
		Dminus[2726] = 14'b0000000_0000000;
		Dminus[2727] = 14'b0000000_0000000;
		Dminus[2728] = 14'b0000000_0000000;
		Dminus[2729] = 14'b0000000_0000000;
		Dminus[2730] = 14'b0000000_0000000;
		Dminus[2731] = 14'b0000000_0000000;
		Dminus[2732] = 14'b0000000_0000000;
		Dminus[2733] = 14'b0000000_0000000;
		Dminus[2734] = 14'b0000000_0000000;
		Dminus[2735] = 14'b0000000_0000000;
		Dminus[2736] = 14'b0000000_0000000;
		Dminus[2737] = 14'b0000000_0000000;
		Dminus[2738] = 14'b0000000_0000000;
		Dminus[2739] = 14'b0000000_0000000;
		Dminus[2740] = 14'b0000000_0000000;
		Dminus[2741] = 14'b0000000_0000000;
		Dminus[2742] = 14'b0000000_0000000;
		Dminus[2743] = 14'b0000000_0000000;
		Dminus[2744] = 14'b0000000_0000000;
		Dminus[2745] = 14'b0000000_0000000;
		Dminus[2746] = 14'b0000000_0000000;
		Dminus[2747] = 14'b0000000_0000000;
		Dminus[2748] = 14'b0000000_0000000;
		Dminus[2749] = 14'b0000000_0000000;
		Dminus[2750] = 14'b0000000_0000000;
		Dminus[2751] = 14'b0000000_0000000;
		Dminus[2752] = 14'b0000000_0000000;
		Dminus[2753] = 14'b0000000_0000000;
		Dminus[2754] = 14'b0000000_0000000;
		Dminus[2755] = 14'b0000000_0000000;
		Dminus[2756] = 14'b0000000_0000000;
		Dminus[2757] = 14'b0000000_0000000;
		Dminus[2758] = 14'b0000000_0000000;
		Dminus[2759] = 14'b0000000_0000000;
		Dminus[2760] = 14'b0000000_0000000;
		Dminus[2761] = 14'b0000000_0000000;
		Dminus[2762] = 14'b0000000_0000000;
		Dminus[2763] = 14'b0000000_0000000;
		Dminus[2764] = 14'b0000000_0000000;
		Dminus[2765] = 14'b0000000_0000000;
		Dminus[2766] = 14'b0000000_0000000;
		Dminus[2767] = 14'b0000000_0000000;
		Dminus[2768] = 14'b0000000_0000000;
		Dminus[2769] = 14'b0000000_0000000;
		Dminus[2770] = 14'b0000000_0000000;
		Dminus[2771] = 14'b0000000_0000000;
		Dminus[2772] = 14'b0000000_0000000;
		Dminus[2773] = 14'b0000000_0000000;
		Dminus[2774] = 14'b0000000_0000000;
		Dminus[2775] = 14'b0000000_0000000;
		Dminus[2776] = 14'b0000000_0000000;
		Dminus[2777] = 14'b0000000_0000000;
		Dminus[2778] = 14'b0000000_0000000;
		Dminus[2779] = 14'b0000000_0000000;
		Dminus[2780] = 14'b0000000_0000000;
		Dminus[2781] = 14'b0000000_0000000;
		Dminus[2782] = 14'b0000000_0000000;
		Dminus[2783] = 14'b0000000_0000000;
		Dminus[2784] = 14'b0000000_0000000;
		Dminus[2785] = 14'b0000000_0000000;
		Dminus[2786] = 14'b0000000_0000000;
		Dminus[2787] = 14'b0000000_0000000;
		Dminus[2788] = 14'b0000000_0000000;
		Dminus[2789] = 14'b0000000_0000000;
		Dminus[2790] = 14'b0000000_0000000;
		Dminus[2791] = 14'b0000000_0000000;
		Dminus[2792] = 14'b0000000_0000000;
		Dminus[2793] = 14'b0000000_0000000;
		Dminus[2794] = 14'b0000000_0000000;
		Dminus[2795] = 14'b0000000_0000000;
		Dminus[2796] = 14'b0000000_0000000;
		Dminus[2797] = 14'b0000000_0000000;
		Dminus[2798] = 14'b0000000_0000000;
		Dminus[2799] = 14'b0000000_0000000;
		Dminus[2800] = 14'b0000000_0000000;
		Dminus[2801] = 14'b0000000_0000000;
		Dminus[2802] = 14'b0000000_0000000;
		Dminus[2803] = 14'b0000000_0000000;
		Dminus[2804] = 14'b0000000_0000000;
		Dminus[2805] = 14'b0000000_0000000;
		Dminus[2806] = 14'b0000000_0000000;
		Dminus[2807] = 14'b0000000_0000000;
		Dminus[2808] = 14'b0000000_0000000;
		Dminus[2809] = 14'b0000000_0000000;
		Dminus[2810] = 14'b0000000_0000000;
		Dminus[2811] = 14'b0000000_0000000;
		Dminus[2812] = 14'b0000000_0000000;
		Dminus[2813] = 14'b0000000_0000000;
		Dminus[2814] = 14'b0000000_0000000;
		Dminus[2815] = 14'b0000000_0000000;
		Dminus[2816] = 14'b0000000_0000000;
		Dminus[2817] = 14'b0000000_0000000;
		Dminus[2818] = 14'b0000000_0000000;
		Dminus[2819] = 14'b0000000_0000000;
		Dminus[2820] = 14'b0000000_0000000;
		Dminus[2821] = 14'b0000000_0000000;
		Dminus[2822] = 14'b0000000_0000000;
		Dminus[2823] = 14'b0000000_0000000;
		Dminus[2824] = 14'b0000000_0000000;
		Dminus[2825] = 14'b0000000_0000000;
		Dminus[2826] = 14'b0000000_0000000;
		Dminus[2827] = 14'b0000000_0000000;
		Dminus[2828] = 14'b0000000_0000000;
		Dminus[2829] = 14'b0000000_0000000;
		Dminus[2830] = 14'b0000000_0000000;
		Dminus[2831] = 14'b0000000_0000000;
		Dminus[2832] = 14'b0000000_0000000;
		Dminus[2833] = 14'b0000000_0000000;
		Dminus[2834] = 14'b0000000_0000000;
		Dminus[2835] = 14'b0000000_0000000;
		Dminus[2836] = 14'b0000000_0000000;
		Dminus[2837] = 14'b0000000_0000000;
		Dminus[2838] = 14'b0000000_0000000;
		Dminus[2839] = 14'b0000000_0000000;
		Dminus[2840] = 14'b0000000_0000000;
		Dminus[2841] = 14'b0000000_0000000;
		Dminus[2842] = 14'b0000000_0000000;
		Dminus[2843] = 14'b0000000_0000000;
		Dminus[2844] = 14'b0000000_0000000;
		Dminus[2845] = 14'b0000000_0000000;
		Dminus[2846] = 14'b0000000_0000000;
		Dminus[2847] = 14'b0000000_0000000;
		Dminus[2848] = 14'b0000000_0000000;
		Dminus[2849] = 14'b0000000_0000000;
		Dminus[2850] = 14'b0000000_0000000;
		Dminus[2851] = 14'b0000000_0000000;
		Dminus[2852] = 14'b0000000_0000000;
		Dminus[2853] = 14'b0000000_0000000;
		Dminus[2854] = 14'b0000000_0000000;
		Dminus[2855] = 14'b0000000_0000000;
		Dminus[2856] = 14'b0000000_0000000;
		Dminus[2857] = 14'b0000000_0000000;
		Dminus[2858] = 14'b0000000_0000000;
		Dminus[2859] = 14'b0000000_0000000;
		Dminus[2860] = 14'b0000000_0000000;
		Dminus[2861] = 14'b0000000_0000000;
		Dminus[2862] = 14'b0000000_0000000;
		Dminus[2863] = 14'b0000000_0000000;
		Dminus[2864] = 14'b0000000_0000000;
		Dminus[2865] = 14'b0000000_0000000;
		Dminus[2866] = 14'b0000000_0000000;
		Dminus[2867] = 14'b0000000_0000000;
		Dminus[2868] = 14'b0000000_0000000;
		Dminus[2869] = 14'b0000000_0000000;
		Dminus[2870] = 14'b0000000_0000000;
		Dminus[2871] = 14'b0000000_0000000;
		Dminus[2872] = 14'b0000000_0000000;
		Dminus[2873] = 14'b0000000_0000000;
		Dminus[2874] = 14'b0000000_0000000;
		Dminus[2875] = 14'b0000000_0000000;
		Dminus[2876] = 14'b0000000_0000000;
		Dminus[2877] = 14'b0000000_0000000;
		Dminus[2878] = 14'b0000000_0000000;
		Dminus[2879] = 14'b0000000_0000000;
		Dminus[2880] = 14'b0000000_0000000;
		Dminus[2881] = 14'b0000000_0000000;
		Dminus[2882] = 14'b0000000_0000000;
		Dminus[2883] = 14'b0000000_0000000;
		Dminus[2884] = 14'b0000000_0000000;
		Dminus[2885] = 14'b0000000_0000000;
		Dminus[2886] = 14'b0000000_0000000;
		Dminus[2887] = 14'b0000000_0000000;
		Dminus[2888] = 14'b0000000_0000000;
		Dminus[2889] = 14'b0000000_0000000;
		Dminus[2890] = 14'b0000000_0000000;
		Dminus[2891] = 14'b0000000_0000000;
		Dminus[2892] = 14'b0000000_0000000;
		Dminus[2893] = 14'b0000000_0000000;
		Dminus[2894] = 14'b0000000_0000000;
		Dminus[2895] = 14'b0000000_0000000;
		Dminus[2896] = 14'b0000000_0000000;
		Dminus[2897] = 14'b0000000_0000000;
		Dminus[2898] = 14'b0000000_0000000;
		Dminus[2899] = 14'b0000000_0000000;
		Dminus[2900] = 14'b0000000_0000000;
		Dminus[2901] = 14'b0000000_0000000;
		Dminus[2902] = 14'b0000000_0000000;
		Dminus[2903] = 14'b0000000_0000000;
		Dminus[2904] = 14'b0000000_0000000;
		Dminus[2905] = 14'b0000000_0000000;
		Dminus[2906] = 14'b0000000_0000000;
		Dminus[2907] = 14'b0000000_0000000;
		Dminus[2908] = 14'b0000000_0000000;
		Dminus[2909] = 14'b0000000_0000000;
		Dminus[2910] = 14'b0000000_0000000;
		Dminus[2911] = 14'b0000000_0000000;
		Dminus[2912] = 14'b0000000_0000000;
		Dminus[2913] = 14'b0000000_0000000;
		Dminus[2914] = 14'b0000000_0000000;
		Dminus[2915] = 14'b0000000_0000000;
		Dminus[2916] = 14'b0000000_0000000;
		Dminus[2917] = 14'b0000000_0000000;
		Dminus[2918] = 14'b0000000_0000000;
		Dminus[2919] = 14'b0000000_0000000;
		Dminus[2920] = 14'b0000000_0000000;
		Dminus[2921] = 14'b0000000_0000000;
		Dminus[2922] = 14'b0000000_0000000;
		Dminus[2923] = 14'b0000000_0000000;
		Dminus[2924] = 14'b0000000_0000000;
		Dminus[2925] = 14'b0000000_0000000;
		Dminus[2926] = 14'b0000000_0000000;
		Dminus[2927] = 14'b0000000_0000000;
		Dminus[2928] = 14'b0000000_0000000;
		Dminus[2929] = 14'b0000000_0000000;
		Dminus[2930] = 14'b0000000_0000000;
		Dminus[2931] = 14'b0000000_0000000;
		Dminus[2932] = 14'b0000000_0000000;
		Dminus[2933] = 14'b0000000_0000000;
		Dminus[2934] = 14'b0000000_0000000;
		Dminus[2935] = 14'b0000000_0000000;
		Dminus[2936] = 14'b0000000_0000000;
		Dminus[2937] = 14'b0000000_0000000;
		Dminus[2938] = 14'b0000000_0000000;
		Dminus[2939] = 14'b0000000_0000000;
		Dminus[2940] = 14'b0000000_0000000;
		Dminus[2941] = 14'b0000000_0000000;
		Dminus[2942] = 14'b0000000_0000000;
		Dminus[2943] = 14'b0000000_0000000;
		Dminus[2944] = 14'b0000000_0000000;
		Dminus[2945] = 14'b0000000_0000000;
		Dminus[2946] = 14'b0000000_0000000;
		Dminus[2947] = 14'b0000000_0000000;
		Dminus[2948] = 14'b0000000_0000000;
		Dminus[2949] = 14'b0000000_0000000;
		Dminus[2950] = 14'b0000000_0000000;
		Dminus[2951] = 14'b0000000_0000000;
		Dminus[2952] = 14'b0000000_0000000;
		Dminus[2953] = 14'b0000000_0000000;
		Dminus[2954] = 14'b0000000_0000000;
		Dminus[2955] = 14'b0000000_0000000;
		Dminus[2956] = 14'b0000000_0000000;
		Dminus[2957] = 14'b0000000_0000000;
		Dminus[2958] = 14'b0000000_0000000;
		Dminus[2959] = 14'b0000000_0000000;
		Dminus[2960] = 14'b0000000_0000000;
		Dminus[2961] = 14'b0000000_0000000;
		Dminus[2962] = 14'b0000000_0000000;
		Dminus[2963] = 14'b0000000_0000000;
		Dminus[2964] = 14'b0000000_0000000;
		Dminus[2965] = 14'b0000000_0000000;
		Dminus[2966] = 14'b0000000_0000000;
		Dminus[2967] = 14'b0000000_0000000;
		Dminus[2968] = 14'b0000000_0000000;
		Dminus[2969] = 14'b0000000_0000000;
		Dminus[2970] = 14'b0000000_0000000;
		Dminus[2971] = 14'b0000000_0000000;
		Dminus[2972] = 14'b0000000_0000000;
		Dminus[2973] = 14'b0000000_0000000;
		Dminus[2974] = 14'b0000000_0000000;
		Dminus[2975] = 14'b0000000_0000000;
		Dminus[2976] = 14'b0000000_0000000;
		Dminus[2977] = 14'b0000000_0000000;
		Dminus[2978] = 14'b0000000_0000000;
		Dminus[2979] = 14'b0000000_0000000;
		Dminus[2980] = 14'b0000000_0000000;
		Dminus[2981] = 14'b0000000_0000000;
		Dminus[2982] = 14'b0000000_0000000;
		Dminus[2983] = 14'b0000000_0000000;
		Dminus[2984] = 14'b0000000_0000000;
		Dminus[2985] = 14'b0000000_0000000;
		Dminus[2986] = 14'b0000000_0000000;
		Dminus[2987] = 14'b0000000_0000000;
		Dminus[2988] = 14'b0000000_0000000;
		Dminus[2989] = 14'b0000000_0000000;
		Dminus[2990] = 14'b0000000_0000000;
		Dminus[2991] = 14'b0000000_0000000;
		Dminus[2992] = 14'b0000000_0000000;
		Dminus[2993] = 14'b0000000_0000000;
		Dminus[2994] = 14'b0000000_0000000;
		Dminus[2995] = 14'b0000000_0000000;
		Dminus[2996] = 14'b0000000_0000000;
		Dminus[2997] = 14'b0000000_0000000;
		Dminus[2998] = 14'b0000000_0000000;
		Dminus[2999] = 14'b0000000_0000000;
		Dminus[3000] = 14'b0000000_0000000;
		Dminus[3001] = 14'b0000000_0000000;
		Dminus[3002] = 14'b0000000_0000000;
		Dminus[3003] = 14'b0000000_0000000;
		Dminus[3004] = 14'b0000000_0000000;
		Dminus[3005] = 14'b0000000_0000000;
		Dminus[3006] = 14'b0000000_0000000;
		Dminus[3007] = 14'b0000000_0000000;
		Dminus[3008] = 14'b0000000_0000000;
		Dminus[3009] = 14'b0000000_0000000;
		Dminus[3010] = 14'b0000000_0000000;
		Dminus[3011] = 14'b0000000_0000000;
		Dminus[3012] = 14'b0000000_0000000;
		Dminus[3013] = 14'b0000000_0000000;
		Dminus[3014] = 14'b0000000_0000000;
		Dminus[3015] = 14'b0000000_0000000;
		Dminus[3016] = 14'b0000000_0000000;
		Dminus[3017] = 14'b0000000_0000000;
		Dminus[3018] = 14'b0000000_0000000;
		Dminus[3019] = 14'b0000000_0000000;
		Dminus[3020] = 14'b0000000_0000000;
		Dminus[3021] = 14'b0000000_0000000;
		Dminus[3022] = 14'b0000000_0000000;
		Dminus[3023] = 14'b0000000_0000000;
		Dminus[3024] = 14'b0000000_0000000;
		Dminus[3025] = 14'b0000000_0000000;
		Dminus[3026] = 14'b0000000_0000000;
		Dminus[3027] = 14'b0000000_0000000;
		Dminus[3028] = 14'b0000000_0000000;
		Dminus[3029] = 14'b0000000_0000000;
		Dminus[3030] = 14'b0000000_0000000;
		Dminus[3031] = 14'b0000000_0000000;
		Dminus[3032] = 14'b0000000_0000000;
		Dminus[3033] = 14'b0000000_0000000;
		Dminus[3034] = 14'b0000000_0000000;
		Dminus[3035] = 14'b0000000_0000000;
		Dminus[3036] = 14'b0000000_0000000;
		Dminus[3037] = 14'b0000000_0000000;
		Dminus[3038] = 14'b0000000_0000000;
		Dminus[3039] = 14'b0000000_0000000;
		Dminus[3040] = 14'b0000000_0000000;
		Dminus[3041] = 14'b0000000_0000000;
		Dminus[3042] = 14'b0000000_0000000;
		Dminus[3043] = 14'b0000000_0000000;
		Dminus[3044] = 14'b0000000_0000000;
		Dminus[3045] = 14'b0000000_0000000;
		Dminus[3046] = 14'b0000000_0000000;
		Dminus[3047] = 14'b0000000_0000000;
		Dminus[3048] = 14'b0000000_0000000;
		Dminus[3049] = 14'b0000000_0000000;
		Dminus[3050] = 14'b0000000_0000000;
		Dminus[3051] = 14'b0000000_0000000;
		Dminus[3052] = 14'b0000000_0000000;
		Dminus[3053] = 14'b0000000_0000000;
		Dminus[3054] = 14'b0000000_0000000;
		Dminus[3055] = 14'b0000000_0000000;
		Dminus[3056] = 14'b0000000_0000000;
		Dminus[3057] = 14'b0000000_0000000;
		Dminus[3058] = 14'b0000000_0000000;
		Dminus[3059] = 14'b0000000_0000000;
		Dminus[3060] = 14'b0000000_0000000;
		Dminus[3061] = 14'b0000000_0000000;
		Dminus[3062] = 14'b0000000_0000000;
		Dminus[3063] = 14'b0000000_0000000;
		Dminus[3064] = 14'b0000000_0000000;
		Dminus[3065] = 14'b0000000_0000000;
		Dminus[3066] = 14'b0000000_0000000;
		Dminus[3067] = 14'b0000000_0000000;
		Dminus[3068] = 14'b0000000_0000000;
		Dminus[3069] = 14'b0000000_0000000;
		Dminus[3070] = 14'b0000000_0000000;
		Dminus[3071] = 14'b0000000_0000000;
		Dminus[3072] = 14'b0000000_0000000;
		Dminus[3073] = 14'b0000000_0000000;
		Dminus[3074] = 14'b0000000_0000000;
		Dminus[3075] = 14'b0000000_0000000;
		Dminus[3076] = 14'b0000000_0000000;
		Dminus[3077] = 14'b0000000_0000000;
		Dminus[3078] = 14'b0000000_0000000;
		Dminus[3079] = 14'b0000000_0000000;
		Dminus[3080] = 14'b0000000_0000000;
		Dminus[3081] = 14'b0000000_0000000;
		Dminus[3082] = 14'b0000000_0000000;
		Dminus[3083] = 14'b0000000_0000000;
		Dminus[3084] = 14'b0000000_0000000;
		Dminus[3085] = 14'b0000000_0000000;
		Dminus[3086] = 14'b0000000_0000000;
		Dminus[3087] = 14'b0000000_0000000;
		Dminus[3088] = 14'b0000000_0000000;
		Dminus[3089] = 14'b0000000_0000000;
		Dminus[3090] = 14'b0000000_0000000;
		Dminus[3091] = 14'b0000000_0000000;
		Dminus[3092] = 14'b0000000_0000000;
		Dminus[3093] = 14'b0000000_0000000;
		Dminus[3094] = 14'b0000000_0000000;
		Dminus[3095] = 14'b0000000_0000000;
		Dminus[3096] = 14'b0000000_0000000;
		Dminus[3097] = 14'b0000000_0000000;
		Dminus[3098] = 14'b0000000_0000000;
		Dminus[3099] = 14'b0000000_0000000;
		Dminus[3100] = 14'b0000000_0000000;
		Dminus[3101] = 14'b0000000_0000000;
		Dminus[3102] = 14'b0000000_0000000;
		Dminus[3103] = 14'b0000000_0000000;
		Dminus[3104] = 14'b0000000_0000000;
		Dminus[3105] = 14'b0000000_0000000;
		Dminus[3106] = 14'b0000000_0000000;
		Dminus[3107] = 14'b0000000_0000000;
		Dminus[3108] = 14'b0000000_0000000;
		Dminus[3109] = 14'b0000000_0000000;
		Dminus[3110] = 14'b0000000_0000000;
		Dminus[3111] = 14'b0000000_0000000;
		Dminus[3112] = 14'b0000000_0000000;
		Dminus[3113] = 14'b0000000_0000000;
		Dminus[3114] = 14'b0000000_0000000;
		Dminus[3115] = 14'b0000000_0000000;
		Dminus[3116] = 14'b0000000_0000000;
		Dminus[3117] = 14'b0000000_0000000;
		Dminus[3118] = 14'b0000000_0000000;
		Dminus[3119] = 14'b0000000_0000000;
		Dminus[3120] = 14'b0000000_0000000;
		Dminus[3121] = 14'b0000000_0000000;
		Dminus[3122] = 14'b0000000_0000000;
		Dminus[3123] = 14'b0000000_0000000;
		Dminus[3124] = 14'b0000000_0000000;
		Dminus[3125] = 14'b0000000_0000000;
		Dminus[3126] = 14'b0000000_0000000;
		Dminus[3127] = 14'b0000000_0000000;
		Dminus[3128] = 14'b0000000_0000000;
		Dminus[3129] = 14'b0000000_0000000;
		Dminus[3130] = 14'b0000000_0000000;
		Dminus[3131] = 14'b0000000_0000000;
		Dminus[3132] = 14'b0000000_0000000;
		Dminus[3133] = 14'b0000000_0000000;
		Dminus[3134] = 14'b0000000_0000000;
		Dminus[3135] = 14'b0000000_0000000;
		Dminus[3136] = 14'b0000000_0000000;
		Dminus[3137] = 14'b0000000_0000000;
		Dminus[3138] = 14'b0000000_0000000;
		Dminus[3139] = 14'b0000000_0000000;
		Dminus[3140] = 14'b0000000_0000000;
		Dminus[3141] = 14'b0000000_0000000;
		Dminus[3142] = 14'b0000000_0000000;
		Dminus[3143] = 14'b0000000_0000000;
		Dminus[3144] = 14'b0000000_0000000;
		Dminus[3145] = 14'b0000000_0000000;
		Dminus[3146] = 14'b0000000_0000000;
		Dminus[3147] = 14'b0000000_0000000;
		Dminus[3148] = 14'b0000000_0000000;
		Dminus[3149] = 14'b0000000_0000000;
		Dminus[3150] = 14'b0000000_0000000;
		Dminus[3151] = 14'b0000000_0000000;
		Dminus[3152] = 14'b0000000_0000000;
		Dminus[3153] = 14'b0000000_0000000;
		Dminus[3154] = 14'b0000000_0000000;
		Dminus[3155] = 14'b0000000_0000000;
		Dminus[3156] = 14'b0000000_0000000;
		Dminus[3157] = 14'b0000000_0000000;
		Dminus[3158] = 14'b0000000_0000000;
		Dminus[3159] = 14'b0000000_0000000;
		Dminus[3160] = 14'b0000000_0000000;
		Dminus[3161] = 14'b0000000_0000000;
		Dminus[3162] = 14'b0000000_0000000;
		Dminus[3163] = 14'b0000000_0000000;
		Dminus[3164] = 14'b0000000_0000000;
		Dminus[3165] = 14'b0000000_0000000;
		Dminus[3166] = 14'b0000000_0000000;
		Dminus[3167] = 14'b0000000_0000000;
		Dminus[3168] = 14'b0000000_0000000;
		Dminus[3169] = 14'b0000000_0000000;
		Dminus[3170] = 14'b0000000_0000000;
		Dminus[3171] = 14'b0000000_0000000;
		Dminus[3172] = 14'b0000000_0000000;
		Dminus[3173] = 14'b0000000_0000000;
		Dminus[3174] = 14'b0000000_0000000;
		Dminus[3175] = 14'b0000000_0000000;
		Dminus[3176] = 14'b0000000_0000000;
		Dminus[3177] = 14'b0000000_0000000;
		Dminus[3178] = 14'b0000000_0000000;
		Dminus[3179] = 14'b0000000_0000000;
		Dminus[3180] = 14'b0000000_0000000;
		Dminus[3181] = 14'b0000000_0000000;
		Dminus[3182] = 14'b0000000_0000000;
		Dminus[3183] = 14'b0000000_0000000;
		Dminus[3184] = 14'b0000000_0000000;
		Dminus[3185] = 14'b0000000_0000000;
		Dminus[3186] = 14'b0000000_0000000;
		Dminus[3187] = 14'b0000000_0000000;
		Dminus[3188] = 14'b0000000_0000000;
		Dminus[3189] = 14'b0000000_0000000;
		Dminus[3190] = 14'b0000000_0000000;
		Dminus[3191] = 14'b0000000_0000000;
		Dminus[3192] = 14'b0000000_0000000;
		Dminus[3193] = 14'b0000000_0000000;
		Dminus[3194] = 14'b0000000_0000000;
		Dminus[3195] = 14'b0000000_0000000;
		Dminus[3196] = 14'b0000000_0000000;
		Dminus[3197] = 14'b0000000_0000000;
		Dminus[3198] = 14'b0000000_0000000;
		Dminus[3199] = 14'b0000000_0000000;
		Dminus[3200] = 14'b0000000_0000000;
		Dminus[3201] = 14'b0000000_0000000;
		Dminus[3202] = 14'b0000000_0000000;
		Dminus[3203] = 14'b0000000_0000000;
		Dminus[3204] = 14'b0000000_0000000;
		Dminus[3205] = 14'b0000000_0000000;
		Dminus[3206] = 14'b0000000_0000000;
		Dminus[3207] = 14'b0000000_0000000;
		Dminus[3208] = 14'b0000000_0000000;
		Dminus[3209] = 14'b0000000_0000000;
		Dminus[3210] = 14'b0000000_0000000;
		Dminus[3211] = 14'b0000000_0000000;
		Dminus[3212] = 14'b0000000_0000000;
		Dminus[3213] = 14'b0000000_0000000;
		Dminus[3214] = 14'b0000000_0000000;
		Dminus[3215] = 14'b0000000_0000000;
		Dminus[3216] = 14'b0000000_0000000;
		Dminus[3217] = 14'b0000000_0000000;
		Dminus[3218] = 14'b0000000_0000000;
		Dminus[3219] = 14'b0000000_0000000;
		Dminus[3220] = 14'b0000000_0000000;
		Dminus[3221] = 14'b0000000_0000000;
		Dminus[3222] = 14'b0000000_0000000;
		Dminus[3223] = 14'b0000000_0000000;
		Dminus[3224] = 14'b0000000_0000000;
		Dminus[3225] = 14'b0000000_0000000;
		Dminus[3226] = 14'b0000000_0000000;
		Dminus[3227] = 14'b0000000_0000000;
		Dminus[3228] = 14'b0000000_0000000;
		Dminus[3229] = 14'b0000000_0000000;
		Dminus[3230] = 14'b0000000_0000000;
		Dminus[3231] = 14'b0000000_0000000;
		Dminus[3232] = 14'b0000000_0000000;
		Dminus[3233] = 14'b0000000_0000000;
		Dminus[3234] = 14'b0000000_0000000;
		Dminus[3235] = 14'b0000000_0000000;
		Dminus[3236] = 14'b0000000_0000000;
		Dminus[3237] = 14'b0000000_0000000;
		Dminus[3238] = 14'b0000000_0000000;
		Dminus[3239] = 14'b0000000_0000000;
		Dminus[3240] = 14'b0000000_0000000;
		Dminus[3241] = 14'b0000000_0000000;
		Dminus[3242] = 14'b0000000_0000000;
		Dminus[3243] = 14'b0000000_0000000;
		Dminus[3244] = 14'b0000000_0000000;
		Dminus[3245] = 14'b0000000_0000000;
		Dminus[3246] = 14'b0000000_0000000;
		Dminus[3247] = 14'b0000000_0000000;
		Dminus[3248] = 14'b0000000_0000000;
		Dminus[3249] = 14'b0000000_0000000;
		Dminus[3250] = 14'b0000000_0000000;
		Dminus[3251] = 14'b0000000_0000000;
		Dminus[3252] = 14'b0000000_0000000;
		Dminus[3253] = 14'b0000000_0000000;
		Dminus[3254] = 14'b0000000_0000000;
		Dminus[3255] = 14'b0000000_0000000;
		Dminus[3256] = 14'b0000000_0000000;
		Dminus[3257] = 14'b0000000_0000000;
		Dminus[3258] = 14'b0000000_0000000;
		Dminus[3259] = 14'b0000000_0000000;
		Dminus[3260] = 14'b0000000_0000000;
		Dminus[3261] = 14'b0000000_0000000;
		Dminus[3262] = 14'b0000000_0000000;
		Dminus[3263] = 14'b0000000_0000000;
		Dminus[3264] = 14'b0000000_0000000;
		Dminus[3265] = 14'b0000000_0000000;
		Dminus[3266] = 14'b0000000_0000000;
		Dminus[3267] = 14'b0000000_0000000;
		Dminus[3268] = 14'b0000000_0000000;
		Dminus[3269] = 14'b0000000_0000000;
		Dminus[3270] = 14'b0000000_0000000;
		Dminus[3271] = 14'b0000000_0000000;
		Dminus[3272] = 14'b0000000_0000000;
		Dminus[3273] = 14'b0000000_0000000;
		Dminus[3274] = 14'b0000000_0000000;
		Dminus[3275] = 14'b0000000_0000000;
		Dminus[3276] = 14'b0000000_0000000;
		Dminus[3277] = 14'b0000000_0000000;
		Dminus[3278] = 14'b0000000_0000000;
		Dminus[3279] = 14'b0000000_0000000;
		Dminus[3280] = 14'b0000000_0000000;
		Dminus[3281] = 14'b0000000_0000000;
		Dminus[3282] = 14'b0000000_0000000;
		Dminus[3283] = 14'b0000000_0000000;
		Dminus[3284] = 14'b0000000_0000000;
		Dminus[3285] = 14'b0000000_0000000;
		Dminus[3286] = 14'b0000000_0000000;
		Dminus[3287] = 14'b0000000_0000000;
		Dminus[3288] = 14'b0000000_0000000;
		Dminus[3289] = 14'b0000000_0000000;
		Dminus[3290] = 14'b0000000_0000000;
		Dminus[3291] = 14'b0000000_0000000;
		Dminus[3292] = 14'b0000000_0000000;
		Dminus[3293] = 14'b0000000_0000000;
		Dminus[3294] = 14'b0000000_0000000;
		Dminus[3295] = 14'b0000000_0000000;
		Dminus[3296] = 14'b0000000_0000000;
		Dminus[3297] = 14'b0000000_0000000;
		Dminus[3298] = 14'b0000000_0000000;
		Dminus[3299] = 14'b0000000_0000000;
		Dminus[3300] = 14'b0000000_0000000;
		Dminus[3301] = 14'b0000000_0000000;
		Dminus[3302] = 14'b0000000_0000000;
		Dminus[3303] = 14'b0000000_0000000;
		Dminus[3304] = 14'b0000000_0000000;
		Dminus[3305] = 14'b0000000_0000000;
		Dminus[3306] = 14'b0000000_0000000;
		Dminus[3307] = 14'b0000000_0000000;
		Dminus[3308] = 14'b0000000_0000000;
		Dminus[3309] = 14'b0000000_0000000;
		Dminus[3310] = 14'b0000000_0000000;
		Dminus[3311] = 14'b0000000_0000000;
		Dminus[3312] = 14'b0000000_0000000;
		Dminus[3313] = 14'b0000000_0000000;
		Dminus[3314] = 14'b0000000_0000000;
		Dminus[3315] = 14'b0000000_0000000;
		Dminus[3316] = 14'b0000000_0000000;
		Dminus[3317] = 14'b0000000_0000000;
		Dminus[3318] = 14'b0000000_0000000;
		Dminus[3319] = 14'b0000000_0000000;
		Dminus[3320] = 14'b0000000_0000000;
		Dminus[3321] = 14'b0000000_0000000;
		Dminus[3322] = 14'b0000000_0000000;
		Dminus[3323] = 14'b0000000_0000000;
		Dminus[3324] = 14'b0000000_0000000;
		Dminus[3325] = 14'b0000000_0000000;
		Dminus[3326] = 14'b0000000_0000000;
		Dminus[3327] = 14'b0000000_0000000;
		Dminus[3328] = 14'b0000000_0000000;
		Dminus[3329] = 14'b0000000_0000000;
		Dminus[3330] = 14'b0000000_0000000;
		Dminus[3331] = 14'b0000000_0000000;
		Dminus[3332] = 14'b0000000_0000000;
		Dminus[3333] = 14'b0000000_0000000;
		Dminus[3334] = 14'b0000000_0000000;
		Dminus[3335] = 14'b0000000_0000000;
		Dminus[3336] = 14'b0000000_0000000;
		Dminus[3337] = 14'b0000000_0000000;
		Dminus[3338] = 14'b0000000_0000000;
		Dminus[3339] = 14'b0000000_0000000;
		Dminus[3340] = 14'b0000000_0000000;
		Dminus[3341] = 14'b0000000_0000000;
		Dminus[3342] = 14'b0000000_0000000;
		Dminus[3343] = 14'b0000000_0000000;
		Dminus[3344] = 14'b0000000_0000000;
		Dminus[3345] = 14'b0000000_0000000;
		Dminus[3346] = 14'b0000000_0000000;
		Dminus[3347] = 14'b0000000_0000000;
		Dminus[3348] = 14'b0000000_0000000;
		Dminus[3349] = 14'b0000000_0000000;
		Dminus[3350] = 14'b0000000_0000000;
		Dminus[3351] = 14'b0000000_0000000;
		Dminus[3352] = 14'b0000000_0000000;
		Dminus[3353] = 14'b0000000_0000000;
		Dminus[3354] = 14'b0000000_0000000;
		Dminus[3355] = 14'b0000000_0000000;
		Dminus[3356] = 14'b0000000_0000000;
		Dminus[3357] = 14'b0000000_0000000;
		Dminus[3358] = 14'b0000000_0000000;
		Dminus[3359] = 14'b0000000_0000000;
		Dminus[3360] = 14'b0000000_0000000;
		Dminus[3361] = 14'b0000000_0000000;
		Dminus[3362] = 14'b0000000_0000000;
		Dminus[3363] = 14'b0000000_0000000;
		Dminus[3364] = 14'b0000000_0000000;
		Dminus[3365] = 14'b0000000_0000000;
		Dminus[3366] = 14'b0000000_0000000;
		Dminus[3367] = 14'b0000000_0000000;
		Dminus[3368] = 14'b0000000_0000000;
		Dminus[3369] = 14'b0000000_0000000;
		Dminus[3370] = 14'b0000000_0000000;
		Dminus[3371] = 14'b0000000_0000000;
		Dminus[3372] = 14'b0000000_0000000;
		Dminus[3373] = 14'b0000000_0000000;
		Dminus[3374] = 14'b0000000_0000000;
		Dminus[3375] = 14'b0000000_0000000;
		Dminus[3376] = 14'b0000000_0000000;
		Dminus[3377] = 14'b0000000_0000000;
		Dminus[3378] = 14'b0000000_0000000;
		Dminus[3379] = 14'b0000000_0000000;
		Dminus[3380] = 14'b0000000_0000000;
		Dminus[3381] = 14'b0000000_0000000;
		Dminus[3382] = 14'b0000000_0000000;
		Dminus[3383] = 14'b0000000_0000000;
		Dminus[3384] = 14'b0000000_0000000;
		Dminus[3385] = 14'b0000000_0000000;
		Dminus[3386] = 14'b0000000_0000000;
		Dminus[3387] = 14'b0000000_0000000;
		Dminus[3388] = 14'b0000000_0000000;
		Dminus[3389] = 14'b0000000_0000000;
		Dminus[3390] = 14'b0000000_0000000;
		Dminus[3391] = 14'b0000000_0000000;
		Dminus[3392] = 14'b0000000_0000000;
		Dminus[3393] = 14'b0000000_0000000;
		Dminus[3394] = 14'b0000000_0000000;
		Dminus[3395] = 14'b0000000_0000000;
		Dminus[3396] = 14'b0000000_0000000;
		Dminus[3397] = 14'b0000000_0000000;
		Dminus[3398] = 14'b0000000_0000000;
		Dminus[3399] = 14'b0000000_0000000;
		Dminus[3400] = 14'b0000000_0000000;
		Dminus[3401] = 14'b0000000_0000000;
		Dminus[3402] = 14'b0000000_0000000;
		Dminus[3403] = 14'b0000000_0000000;
		Dminus[3404] = 14'b0000000_0000000;
		Dminus[3405] = 14'b0000000_0000000;
		Dminus[3406] = 14'b0000000_0000000;
		Dminus[3407] = 14'b0000000_0000000;
		Dminus[3408] = 14'b0000000_0000000;
		Dminus[3409] = 14'b0000000_0000000;
		Dminus[3410] = 14'b0000000_0000000;
		Dminus[3411] = 14'b0000000_0000000;
		Dminus[3412] = 14'b0000000_0000000;
		Dminus[3413] = 14'b0000000_0000000;
		Dminus[3414] = 14'b0000000_0000000;
		Dminus[3415] = 14'b0000000_0000000;
		Dminus[3416] = 14'b0000000_0000000;
		Dminus[3417] = 14'b0000000_0000000;
		Dminus[3418] = 14'b0000000_0000000;
		Dminus[3419] = 14'b0000000_0000000;
		Dminus[3420] = 14'b0000000_0000000;
		Dminus[3421] = 14'b0000000_0000000;
		Dminus[3422] = 14'b0000000_0000000;
		Dminus[3423] = 14'b0000000_0000000;
		Dminus[3424] = 14'b0000000_0000000;
		Dminus[3425] = 14'b0000000_0000000;
		Dminus[3426] = 14'b0000000_0000000;
		Dminus[3427] = 14'b0000000_0000000;
		Dminus[3428] = 14'b0000000_0000000;
		Dminus[3429] = 14'b0000000_0000000;
		Dminus[3430] = 14'b0000000_0000000;
		Dminus[3431] = 14'b0000000_0000000;
		Dminus[3432] = 14'b0000000_0000000;
		Dminus[3433] = 14'b0000000_0000000;
		Dminus[3434] = 14'b0000000_0000000;
		Dminus[3435] = 14'b0000000_0000000;
		Dminus[3436] = 14'b0000000_0000000;
		Dminus[3437] = 14'b0000000_0000000;
		Dminus[3438] = 14'b0000000_0000000;
		Dminus[3439] = 14'b0000000_0000000;
		Dminus[3440] = 14'b0000000_0000000;
		Dminus[3441] = 14'b0000000_0000000;
		Dminus[3442] = 14'b0000000_0000000;
		Dminus[3443] = 14'b0000000_0000000;
		Dminus[3444] = 14'b0000000_0000000;
		Dminus[3445] = 14'b0000000_0000000;
		Dminus[3446] = 14'b0000000_0000000;
		Dminus[3447] = 14'b0000000_0000000;
		Dminus[3448] = 14'b0000000_0000000;
		Dminus[3449] = 14'b0000000_0000000;
		Dminus[3450] = 14'b0000000_0000000;
		Dminus[3451] = 14'b0000000_0000000;
		Dminus[3452] = 14'b0000000_0000000;
		Dminus[3453] = 14'b0000000_0000000;
		Dminus[3454] = 14'b0000000_0000000;
		Dminus[3455] = 14'b0000000_0000000;
		Dminus[3456] = 14'b0000000_0000000;
		Dminus[3457] = 14'b0000000_0000000;
		Dminus[3458] = 14'b0000000_0000000;
		Dminus[3459] = 14'b0000000_0000000;
		Dminus[3460] = 14'b0000000_0000000;
		Dminus[3461] = 14'b0000000_0000000;
		Dminus[3462] = 14'b0000000_0000000;
		Dminus[3463] = 14'b0000000_0000000;
		Dminus[3464] = 14'b0000000_0000000;
		Dminus[3465] = 14'b0000000_0000000;
		Dminus[3466] = 14'b0000000_0000000;
		Dminus[3467] = 14'b0000000_0000000;
		Dminus[3468] = 14'b0000000_0000000;
		Dminus[3469] = 14'b0000000_0000000;
		Dminus[3470] = 14'b0000000_0000000;
		Dminus[3471] = 14'b0000000_0000000;
		Dminus[3472] = 14'b0000000_0000000;
		Dminus[3473] = 14'b0000000_0000000;
		Dminus[3474] = 14'b0000000_0000000;
		Dminus[3475] = 14'b0000000_0000000;
		Dminus[3476] = 14'b0000000_0000000;
		Dminus[3477] = 14'b0000000_0000000;
		Dminus[3478] = 14'b0000000_0000000;
		Dminus[3479] = 14'b0000000_0000000;
		Dminus[3480] = 14'b0000000_0000000;
		Dminus[3481] = 14'b0000000_0000000;
		Dminus[3482] = 14'b0000000_0000000;
		Dminus[3483] = 14'b0000000_0000000;
		Dminus[3484] = 14'b0000000_0000000;
		Dminus[3485] = 14'b0000000_0000000;
		Dminus[3486] = 14'b0000000_0000000;
		Dminus[3487] = 14'b0000000_0000000;
		Dminus[3488] = 14'b0000000_0000000;
		Dminus[3489] = 14'b0000000_0000000;
		Dminus[3490] = 14'b0000000_0000000;
		Dminus[3491] = 14'b0000000_0000000;
		Dminus[3492] = 14'b0000000_0000000;
		Dminus[3493] = 14'b0000000_0000000;
		Dminus[3494] = 14'b0000000_0000000;
		Dminus[3495] = 14'b0000000_0000000;
		Dminus[3496] = 14'b0000000_0000000;
		Dminus[3497] = 14'b0000000_0000000;
		Dminus[3498] = 14'b0000000_0000000;
		Dminus[3499] = 14'b0000000_0000000;
		Dminus[3500] = 14'b0000000_0000000;
		Dminus[3501] = 14'b0000000_0000000;
		Dminus[3502] = 14'b0000000_0000000;
		Dminus[3503] = 14'b0000000_0000000;
		Dminus[3504] = 14'b0000000_0000000;
		Dminus[3505] = 14'b0000000_0000000;
		Dminus[3506] = 14'b0000000_0000000;
		Dminus[3507] = 14'b0000000_0000000;
		Dminus[3508] = 14'b0000000_0000000;
		Dminus[3509] = 14'b0000000_0000000;
		Dminus[3510] = 14'b0000000_0000000;
		Dminus[3511] = 14'b0000000_0000000;
		Dminus[3512] = 14'b0000000_0000000;
		Dminus[3513] = 14'b0000000_0000000;
		Dminus[3514] = 14'b0000000_0000000;
		Dminus[3515] = 14'b0000000_0000000;
		Dminus[3516] = 14'b0000000_0000000;
		Dminus[3517] = 14'b0000000_0000000;
		Dminus[3518] = 14'b0000000_0000000;
		Dminus[3519] = 14'b0000000_0000000;
		Dminus[3520] = 14'b0000000_0000000;
		Dminus[3521] = 14'b0000000_0000000;
		Dminus[3522] = 14'b0000000_0000000;
		Dminus[3523] = 14'b0000000_0000000;
		Dminus[3524] = 14'b0000000_0000000;
		Dminus[3525] = 14'b0000000_0000000;
		Dminus[3526] = 14'b0000000_0000000;
		Dminus[3527] = 14'b0000000_0000000;
		Dminus[3528] = 14'b0000000_0000000;
		Dminus[3529] = 14'b0000000_0000000;
		Dminus[3530] = 14'b0000000_0000000;
		Dminus[3531] = 14'b0000000_0000000;
		Dminus[3532] = 14'b0000000_0000000;
		Dminus[3533] = 14'b0000000_0000000;
		Dminus[3534] = 14'b0000000_0000000;
		Dminus[3535] = 14'b0000000_0000000;
		Dminus[3536] = 14'b0000000_0000000;
		Dminus[3537] = 14'b0000000_0000000;
		Dminus[3538] = 14'b0000000_0000000;
		Dminus[3539] = 14'b0000000_0000000;
		Dminus[3540] = 14'b0000000_0000000;
		Dminus[3541] = 14'b0000000_0000000;
		Dminus[3542] = 14'b0000000_0000000;
		Dminus[3543] = 14'b0000000_0000000;
		Dminus[3544] = 14'b0000000_0000000;
		Dminus[3545] = 14'b0000000_0000000;
		Dminus[3546] = 14'b0000000_0000000;
		Dminus[3547] = 14'b0000000_0000000;
		Dminus[3548] = 14'b0000000_0000000;
		Dminus[3549] = 14'b0000000_0000000;
		Dminus[3550] = 14'b0000000_0000000;
		Dminus[3551] = 14'b0000000_0000000;
		Dminus[3552] = 14'b0000000_0000000;
		Dminus[3553] = 14'b0000000_0000000;
		Dminus[3554] = 14'b0000000_0000000;
		Dminus[3555] = 14'b0000000_0000000;
		Dminus[3556] = 14'b0000000_0000000;
		Dminus[3557] = 14'b0000000_0000000;
		Dminus[3558] = 14'b0000000_0000000;
		Dminus[3559] = 14'b0000000_0000000;
		Dminus[3560] = 14'b0000000_0000000;
		Dminus[3561] = 14'b0000000_0000000;
		Dminus[3562] = 14'b0000000_0000000;
		Dminus[3563] = 14'b0000000_0000000;
		Dminus[3564] = 14'b0000000_0000000;
		Dminus[3565] = 14'b0000000_0000000;
		Dminus[3566] = 14'b0000000_0000000;
		Dminus[3567] = 14'b0000000_0000000;
		Dminus[3568] = 14'b0000000_0000000;
		Dminus[3569] = 14'b0000000_0000000;
		Dminus[3570] = 14'b0000000_0000000;
		Dminus[3571] = 14'b0000000_0000000;
		Dminus[3572] = 14'b0000000_0000000;
		Dminus[3573] = 14'b0000000_0000000;
		Dminus[3574] = 14'b0000000_0000000;
		Dminus[3575] = 14'b0000000_0000000;
		Dminus[3576] = 14'b0000000_0000000;
		Dminus[3577] = 14'b0000000_0000000;
		Dminus[3578] = 14'b0000000_0000000;
		Dminus[3579] = 14'b0000000_0000000;
		Dminus[3580] = 14'b0000000_0000000;
		Dminus[3581] = 14'b0000000_0000000;
		Dminus[3582] = 14'b0000000_0000000;
		Dminus[3583] = 14'b0000000_0000000;
		Dminus[3584] = 14'b0000000_0000000;
		Dminus[3585] = 14'b0000000_0000000;
		Dminus[3586] = 14'b0000000_0000000;
		Dminus[3587] = 14'b0000000_0000000;
		Dminus[3588] = 14'b0000000_0000000;
		Dminus[3589] = 14'b0000000_0000000;
		Dminus[3590] = 14'b0000000_0000000;
		Dminus[3591] = 14'b0000000_0000000;
		Dminus[3592] = 14'b0000000_0000000;
		Dminus[3593] = 14'b0000000_0000000;
		Dminus[3594] = 14'b0000000_0000000;
		Dminus[3595] = 14'b0000000_0000000;
		Dminus[3596] = 14'b0000000_0000000;
		Dminus[3597] = 14'b0000000_0000000;
		Dminus[3598] = 14'b0000000_0000000;
		Dminus[3599] = 14'b0000000_0000000;
		Dminus[3600] = 14'b0000000_0000000;
		Dminus[3601] = 14'b0000000_0000000;
		Dminus[3602] = 14'b0000000_0000000;
		Dminus[3603] = 14'b0000000_0000000;
		Dminus[3604] = 14'b0000000_0000000;
		Dminus[3605] = 14'b0000000_0000000;
		Dminus[3606] = 14'b0000000_0000000;
		Dminus[3607] = 14'b0000000_0000000;
		Dminus[3608] = 14'b0000000_0000000;
		Dminus[3609] = 14'b0000000_0000000;
		Dminus[3610] = 14'b0000000_0000000;
		Dminus[3611] = 14'b0000000_0000000;
		Dminus[3612] = 14'b0000000_0000000;
		Dminus[3613] = 14'b0000000_0000000;
		Dminus[3614] = 14'b0000000_0000000;
		Dminus[3615] = 14'b0000000_0000000;
		Dminus[3616] = 14'b0000000_0000000;
		Dminus[3617] = 14'b0000000_0000000;
		Dminus[3618] = 14'b0000000_0000000;
		Dminus[3619] = 14'b0000000_0000000;
		Dminus[3620] = 14'b0000000_0000000;
		Dminus[3621] = 14'b0000000_0000000;
		Dminus[3622] = 14'b0000000_0000000;
		Dminus[3623] = 14'b0000000_0000000;
		Dminus[3624] = 14'b0000000_0000000;
		Dminus[3625] = 14'b0000000_0000000;
		Dminus[3626] = 14'b0000000_0000000;
		Dminus[3627] = 14'b0000000_0000000;
		Dminus[3628] = 14'b0000000_0000000;
		Dminus[3629] = 14'b0000000_0000000;
		Dminus[3630] = 14'b0000000_0000000;
		Dminus[3631] = 14'b0000000_0000000;
		Dminus[3632] = 14'b0000000_0000000;
		Dminus[3633] = 14'b0000000_0000000;
		Dminus[3634] = 14'b0000000_0000000;
		Dminus[3635] = 14'b0000000_0000000;
		Dminus[3636] = 14'b0000000_0000000;
		Dminus[3637] = 14'b0000000_0000000;
		Dminus[3638] = 14'b0000000_0000000;
		Dminus[3639] = 14'b0000000_0000000;
		Dminus[3640] = 14'b0000000_0000000;
		Dminus[3641] = 14'b0000000_0000000;
		Dminus[3642] = 14'b0000000_0000000;
		Dminus[3643] = 14'b0000000_0000000;
		Dminus[3644] = 14'b0000000_0000000;
		Dminus[3645] = 14'b0000000_0000000;
		Dminus[3646] = 14'b0000000_0000000;
		Dminus[3647] = 14'b0000000_0000000;
		Dminus[3648] = 14'b0000000_0000000;
		Dminus[3649] = 14'b0000000_0000000;
		Dminus[3650] = 14'b0000000_0000000;
		Dminus[3651] = 14'b0000000_0000000;
		Dminus[3652] = 14'b0000000_0000000;
		Dminus[3653] = 14'b0000000_0000000;
		Dminus[3654] = 14'b0000000_0000000;
		Dminus[3655] = 14'b0000000_0000000;
		Dminus[3656] = 14'b0000000_0000000;
		Dminus[3657] = 14'b0000000_0000000;
		Dminus[3658] = 14'b0000000_0000000;
		Dminus[3659] = 14'b0000000_0000000;
		Dminus[3660] = 14'b0000000_0000000;
		Dminus[3661] = 14'b0000000_0000000;
		Dminus[3662] = 14'b0000000_0000000;
		Dminus[3663] = 14'b0000000_0000000;
		Dminus[3664] = 14'b0000000_0000000;
		Dminus[3665] = 14'b0000000_0000000;
		Dminus[3666] = 14'b0000000_0000000;
		Dminus[3667] = 14'b0000000_0000000;
		Dminus[3668] = 14'b0000000_0000000;
		Dminus[3669] = 14'b0000000_0000000;
		Dminus[3670] = 14'b0000000_0000000;
		Dminus[3671] = 14'b0000000_0000000;
		Dminus[3672] = 14'b0000000_0000000;
		Dminus[3673] = 14'b0000000_0000000;
		Dminus[3674] = 14'b0000000_0000000;
		Dminus[3675] = 14'b0000000_0000000;
		Dminus[3676] = 14'b0000000_0000000;
		Dminus[3677] = 14'b0000000_0000000;
		Dminus[3678] = 14'b0000000_0000000;
		Dminus[3679] = 14'b0000000_0000000;
		Dminus[3680] = 14'b0000000_0000000;
		Dminus[3681] = 14'b0000000_0000000;
		Dminus[3682] = 14'b0000000_0000000;
		Dminus[3683] = 14'b0000000_0000000;
		Dminus[3684] = 14'b0000000_0000000;
		Dminus[3685] = 14'b0000000_0000000;
		Dminus[3686] = 14'b0000000_0000000;
		Dminus[3687] = 14'b0000000_0000000;
		Dminus[3688] = 14'b0000000_0000000;
		Dminus[3689] = 14'b0000000_0000000;
		Dminus[3690] = 14'b0000000_0000000;
		Dminus[3691] = 14'b0000000_0000000;
		Dminus[3692] = 14'b0000000_0000000;
		Dminus[3693] = 14'b0000000_0000000;
		Dminus[3694] = 14'b0000000_0000000;
		Dminus[3695] = 14'b0000000_0000000;
		Dminus[3696] = 14'b0000000_0000000;
		Dminus[3697] = 14'b0000000_0000000;
		Dminus[3698] = 14'b0000000_0000000;
		Dminus[3699] = 14'b0000000_0000000;
		Dminus[3700] = 14'b0000000_0000000;
		Dminus[3701] = 14'b0000000_0000000;
		Dminus[3702] = 14'b0000000_0000000;
		Dminus[3703] = 14'b0000000_0000000;
		Dminus[3704] = 14'b0000000_0000000;
		Dminus[3705] = 14'b0000000_0000000;
		Dminus[3706] = 14'b0000000_0000000;
		Dminus[3707] = 14'b0000000_0000000;
		Dminus[3708] = 14'b0000000_0000000;
		Dminus[3709] = 14'b0000000_0000000;
		Dminus[3710] = 14'b0000000_0000000;
		Dminus[3711] = 14'b0000000_0000000;
		Dminus[3712] = 14'b0000000_0000000;
		Dminus[3713] = 14'b0000000_0000000;
		Dminus[3714] = 14'b0000000_0000000;
		Dminus[3715] = 14'b0000000_0000000;
		Dminus[3716] = 14'b0000000_0000000;
		Dminus[3717] = 14'b0000000_0000000;
		Dminus[3718] = 14'b0000000_0000000;
		Dminus[3719] = 14'b0000000_0000000;
		Dminus[3720] = 14'b0000000_0000000;
		Dminus[3721] = 14'b0000000_0000000;
		Dminus[3722] = 14'b0000000_0000000;
		Dminus[3723] = 14'b0000000_0000000;
		Dminus[3724] = 14'b0000000_0000000;
		Dminus[3725] = 14'b0000000_0000000;
		Dminus[3726] = 14'b0000000_0000000;
		Dminus[3727] = 14'b0000000_0000000;
		Dminus[3728] = 14'b0000000_0000000;
		Dminus[3729] = 14'b0000000_0000000;
		Dminus[3730] = 14'b0000000_0000000;
		Dminus[3731] = 14'b0000000_0000000;
		Dminus[3732] = 14'b0000000_0000000;
		Dminus[3733] = 14'b0000000_0000000;
		Dminus[3734] = 14'b0000000_0000000;
		Dminus[3735] = 14'b0000000_0000000;
		Dminus[3736] = 14'b0000000_0000000;
		Dminus[3737] = 14'b0000000_0000000;
		Dminus[3738] = 14'b0000000_0000000;
		Dminus[3739] = 14'b0000000_0000000;
		Dminus[3740] = 14'b0000000_0000000;
		Dminus[3741] = 14'b0000000_0000000;
		Dminus[3742] = 14'b0000000_0000000;
		Dminus[3743] = 14'b0000000_0000000;
		Dminus[3744] = 14'b0000000_0000000;
		Dminus[3745] = 14'b0000000_0000000;
		Dminus[3746] = 14'b0000000_0000000;
		Dminus[3747] = 14'b0000000_0000000;
		Dminus[3748] = 14'b0000000_0000000;
		Dminus[3749] = 14'b0000000_0000000;
		Dminus[3750] = 14'b0000000_0000000;
		Dminus[3751] = 14'b0000000_0000000;
		Dminus[3752] = 14'b0000000_0000000;
		Dminus[3753] = 14'b0000000_0000000;
		Dminus[3754] = 14'b0000000_0000000;
		Dminus[3755] = 14'b0000000_0000000;
		Dminus[3756] = 14'b0000000_0000000;
		Dminus[3757] = 14'b0000000_0000000;
		Dminus[3758] = 14'b0000000_0000000;
		Dminus[3759] = 14'b0000000_0000000;
		Dminus[3760] = 14'b0000000_0000000;
		Dminus[3761] = 14'b0000000_0000000;
		Dminus[3762] = 14'b0000000_0000000;
		Dminus[3763] = 14'b0000000_0000000;
		Dminus[3764] = 14'b0000000_0000000;
		Dminus[3765] = 14'b0000000_0000000;
		Dminus[3766] = 14'b0000000_0000000;
		Dminus[3767] = 14'b0000000_0000000;
		Dminus[3768] = 14'b0000000_0000000;
		Dminus[3769] = 14'b0000000_0000000;
		Dminus[3770] = 14'b0000000_0000000;
		Dminus[3771] = 14'b0000000_0000000;
		Dminus[3772] = 14'b0000000_0000000;
		Dminus[3773] = 14'b0000000_0000000;
		Dminus[3774] = 14'b0000000_0000000;
		Dminus[3775] = 14'b0000000_0000000;
		Dminus[3776] = 14'b0000000_0000000;
		Dminus[3777] = 14'b0000000_0000000;
		Dminus[3778] = 14'b0000000_0000000;
		Dminus[3779] = 14'b0000000_0000000;
		Dminus[3780] = 14'b0000000_0000000;
		Dminus[3781] = 14'b0000000_0000000;
		Dminus[3782] = 14'b0000000_0000000;
		Dminus[3783] = 14'b0000000_0000000;
		Dminus[3784] = 14'b0000000_0000000;
		Dminus[3785] = 14'b0000000_0000000;
		Dminus[3786] = 14'b0000000_0000000;
		Dminus[3787] = 14'b0000000_0000000;
		Dminus[3788] = 14'b0000000_0000000;
		Dminus[3789] = 14'b0000000_0000000;
		Dminus[3790] = 14'b0000000_0000000;
		Dminus[3791] = 14'b0000000_0000000;
		Dminus[3792] = 14'b0000000_0000000;
		Dminus[3793] = 14'b0000000_0000000;
		Dminus[3794] = 14'b0000000_0000000;
		Dminus[3795] = 14'b0000000_0000000;
		Dminus[3796] = 14'b0000000_0000000;
		Dminus[3797] = 14'b0000000_0000000;
		Dminus[3798] = 14'b0000000_0000000;
		Dminus[3799] = 14'b0000000_0000000;
		Dminus[3800] = 14'b0000000_0000000;
		Dminus[3801] = 14'b0000000_0000000;
		Dminus[3802] = 14'b0000000_0000000;
		Dminus[3803] = 14'b0000000_0000000;
		Dminus[3804] = 14'b0000000_0000000;
		Dminus[3805] = 14'b0000000_0000000;
		Dminus[3806] = 14'b0000000_0000000;
		Dminus[3807] = 14'b0000000_0000000;
		Dminus[3808] = 14'b0000000_0000000;
		Dminus[3809] = 14'b0000000_0000000;
		Dminus[3810] = 14'b0000000_0000000;
		Dminus[3811] = 14'b0000000_0000000;
		Dminus[3812] = 14'b0000000_0000000;
		Dminus[3813] = 14'b0000000_0000000;
		Dminus[3814] = 14'b0000000_0000000;
		Dminus[3815] = 14'b0000000_0000000;
		Dminus[3816] = 14'b0000000_0000000;
		Dminus[3817] = 14'b0000000_0000000;
		Dminus[3818] = 14'b0000000_0000000;
		Dminus[3819] = 14'b0000000_0000000;
		Dminus[3820] = 14'b0000000_0000000;
		Dminus[3821] = 14'b0000000_0000000;
		Dminus[3822] = 14'b0000000_0000000;
		Dminus[3823] = 14'b0000000_0000000;
		Dminus[3824] = 14'b0000000_0000000;
		Dminus[3825] = 14'b0000000_0000000;
		Dminus[3826] = 14'b0000000_0000000;
		Dminus[3827] = 14'b0000000_0000000;
		Dminus[3828] = 14'b0000000_0000000;
		Dminus[3829] = 14'b0000000_0000000;
		Dminus[3830] = 14'b0000000_0000000;
		Dminus[3831] = 14'b0000000_0000000;
		Dminus[3832] = 14'b0000000_0000000;
		Dminus[3833] = 14'b0000000_0000000;
		Dminus[3834] = 14'b0000000_0000000;
		Dminus[3835] = 14'b0000000_0000000;
		Dminus[3836] = 14'b0000000_0000000;
		Dminus[3837] = 14'b0000000_0000000;
		Dminus[3838] = 14'b0000000_0000000;
		Dminus[3839] = 14'b0000000_0000000;
		Dminus[3840] = 14'b0000000_0000000;
		Dminus[3841] = 14'b0000000_0000000;
		Dminus[3842] = 14'b0000000_0000000;
		Dminus[3843] = 14'b0000000_0000000;
		Dminus[3844] = 14'b0000000_0000000;
		Dminus[3845] = 14'b0000000_0000000;
		Dminus[3846] = 14'b0000000_0000000;
		Dminus[3847] = 14'b0000000_0000000;
		Dminus[3848] = 14'b0000000_0000000;
		Dminus[3849] = 14'b0000000_0000000;
		Dminus[3850] = 14'b0000000_0000000;
		Dminus[3851] = 14'b0000000_0000000;
		Dminus[3852] = 14'b0000000_0000000;
		Dminus[3853] = 14'b0000000_0000000;
		Dminus[3854] = 14'b0000000_0000000;
		Dminus[3855] = 14'b0000000_0000000;
		Dminus[3856] = 14'b0000000_0000000;
		Dminus[3857] = 14'b0000000_0000000;
		Dminus[3858] = 14'b0000000_0000000;
		Dminus[3859] = 14'b0000000_0000000;
		Dminus[3860] = 14'b0000000_0000000;
		Dminus[3861] = 14'b0000000_0000000;
		Dminus[3862] = 14'b0000000_0000000;
		Dminus[3863] = 14'b0000000_0000000;
		Dminus[3864] = 14'b0000000_0000000;
		Dminus[3865] = 14'b0000000_0000000;
		Dminus[3866] = 14'b0000000_0000000;
		Dminus[3867] = 14'b0000000_0000000;
		Dminus[3868] = 14'b0000000_0000000;
		Dminus[3869] = 14'b0000000_0000000;
		Dminus[3870] = 14'b0000000_0000000;
		Dminus[3871] = 14'b0000000_0000000;
		Dminus[3872] = 14'b0000000_0000000;
		Dminus[3873] = 14'b0000000_0000000;
		Dminus[3874] = 14'b0000000_0000000;
		Dminus[3875] = 14'b0000000_0000000;
		Dminus[3876] = 14'b0000000_0000000;
		Dminus[3877] = 14'b0000000_0000000;
		Dminus[3878] = 14'b0000000_0000000;
		Dminus[3879] = 14'b0000000_0000000;
		Dminus[3880] = 14'b0000000_0000000;
		Dminus[3881] = 14'b0000000_0000000;
		Dminus[3882] = 14'b0000000_0000000;
		Dminus[3883] = 14'b0000000_0000000;
		Dminus[3884] = 14'b0000000_0000000;
		Dminus[3885] = 14'b0000000_0000000;
		Dminus[3886] = 14'b0000000_0000000;
		Dminus[3887] = 14'b0000000_0000000;
		Dminus[3888] = 14'b0000000_0000000;
		Dminus[3889] = 14'b0000000_0000000;
		Dminus[3890] = 14'b0000000_0000000;
		Dminus[3891] = 14'b0000000_0000000;
		Dminus[3892] = 14'b0000000_0000000;
		Dminus[3893] = 14'b0000000_0000000;
		Dminus[3894] = 14'b0000000_0000000;
		Dminus[3895] = 14'b0000000_0000000;
		Dminus[3896] = 14'b0000000_0000000;
		Dminus[3897] = 14'b0000000_0000000;
		Dminus[3898] = 14'b0000000_0000000;
		Dminus[3899] = 14'b0000000_0000000;
		Dminus[3900] = 14'b0000000_0000000;
		Dminus[3901] = 14'b0000000_0000000;
		Dminus[3902] = 14'b0000000_0000000;
		Dminus[3903] = 14'b0000000_0000000;
		Dminus[3904] = 14'b0000000_0000000;
		Dminus[3905] = 14'b0000000_0000000;
		Dminus[3906] = 14'b0000000_0000000;
		Dminus[3907] = 14'b0000000_0000000;
		Dminus[3908] = 14'b0000000_0000000;
		Dminus[3909] = 14'b0000000_0000000;
		Dminus[3910] = 14'b0000000_0000000;
		Dminus[3911] = 14'b0000000_0000000;
		Dminus[3912] = 14'b0000000_0000000;
		Dminus[3913] = 14'b0000000_0000000;
		Dminus[3914] = 14'b0000000_0000000;
		Dminus[3915] = 14'b0000000_0000000;
		Dminus[3916] = 14'b0000000_0000000;
		Dminus[3917] = 14'b0000000_0000000;
		Dminus[3918] = 14'b0000000_0000000;
		Dminus[3919] = 14'b0000000_0000000;
		Dminus[3920] = 14'b0000000_0000000;
		Dminus[3921] = 14'b0000000_0000000;
		Dminus[3922] = 14'b0000000_0000000;
		Dminus[3923] = 14'b0000000_0000000;
		Dminus[3924] = 14'b0000000_0000000;
		Dminus[3925] = 14'b0000000_0000000;
		Dminus[3926] = 14'b0000000_0000000;
		Dminus[3927] = 14'b0000000_0000000;
		Dminus[3928] = 14'b0000000_0000000;
		Dminus[3929] = 14'b0000000_0000000;
		Dminus[3930] = 14'b0000000_0000000;
		Dminus[3931] = 14'b0000000_0000000;
		Dminus[3932] = 14'b0000000_0000000;
		Dminus[3933] = 14'b0000000_0000000;
		Dminus[3934] = 14'b0000000_0000000;
		Dminus[3935] = 14'b0000000_0000000;
		Dminus[3936] = 14'b0000000_0000000;
		Dminus[3937] = 14'b0000000_0000000;
		Dminus[3938] = 14'b0000000_0000000;
		Dminus[3939] = 14'b0000000_0000000;
		Dminus[3940] = 14'b0000000_0000000;
		Dminus[3941] = 14'b0000000_0000000;
		Dminus[3942] = 14'b0000000_0000000;
		Dminus[3943] = 14'b0000000_0000000;
		Dminus[3944] = 14'b0000000_0000000;
		Dminus[3945] = 14'b0000000_0000000;
		Dminus[3946] = 14'b0000000_0000000;
		Dminus[3947] = 14'b0000000_0000000;
		Dminus[3948] = 14'b0000000_0000000;
		Dminus[3949] = 14'b0000000_0000000;
		Dminus[3950] = 14'b0000000_0000000;
		Dminus[3951] = 14'b0000000_0000000;
		Dminus[3952] = 14'b0000000_0000000;
		Dminus[3953] = 14'b0000000_0000000;
		Dminus[3954] = 14'b0000000_0000000;
		Dminus[3955] = 14'b0000000_0000000;
		Dminus[3956] = 14'b0000000_0000000;
		Dminus[3957] = 14'b0000000_0000000;
		Dminus[3958] = 14'b0000000_0000000;
		Dminus[3959] = 14'b0000000_0000000;
		Dminus[3960] = 14'b0000000_0000000;
		Dminus[3961] = 14'b0000000_0000000;
		Dminus[3962] = 14'b0000000_0000000;
		Dminus[3963] = 14'b0000000_0000000;
		Dminus[3964] = 14'b0000000_0000000;
		Dminus[3965] = 14'b0000000_0000000;
		Dminus[3966] = 14'b0000000_0000000;
		Dminus[3967] = 14'b0000000_0000000;
		Dminus[3968] = 14'b0000000_0000000;
		Dminus[3969] = 14'b0000000_0000000;
		Dminus[3970] = 14'b0000000_0000000;
		Dminus[3971] = 14'b0000000_0000000;
		Dminus[3972] = 14'b0000000_0000000;
		Dminus[3973] = 14'b0000000_0000000;
		Dminus[3974] = 14'b0000000_0000000;
		Dminus[3975] = 14'b0000000_0000000;
		Dminus[3976] = 14'b0000000_0000000;
		Dminus[3977] = 14'b0000000_0000000;
		Dminus[3978] = 14'b0000000_0000000;
		Dminus[3979] = 14'b0000000_0000000;
		Dminus[3980] = 14'b0000000_0000000;
		Dminus[3981] = 14'b0000000_0000000;
		Dminus[3982] = 14'b0000000_0000000;
		Dminus[3983] = 14'b0000000_0000000;
		Dminus[3984] = 14'b0000000_0000000;
		Dminus[3985] = 14'b0000000_0000000;
		Dminus[3986] = 14'b0000000_0000000;
		Dminus[3987] = 14'b0000000_0000000;
		Dminus[3988] = 14'b0000000_0000000;
		Dminus[3989] = 14'b0000000_0000000;
		Dminus[3990] = 14'b0000000_0000000;
		Dminus[3991] = 14'b0000000_0000000;
		Dminus[3992] = 14'b0000000_0000000;
		Dminus[3993] = 14'b0000000_0000000;
		Dminus[3994] = 14'b0000000_0000000;
		Dminus[3995] = 14'b0000000_0000000;
		Dminus[3996] = 14'b0000000_0000000;
		Dminus[3997] = 14'b0000000_0000000;
		Dminus[3998] = 14'b0000000_0000000;
		Dminus[3999] = 14'b0000000_0000000;
		Dminus[4000] = 14'b0000000_0000000;
		Dminus[4001] = 14'b0000000_0000000;
		Dminus[4002] = 14'b0000000_0000000;
		Dminus[4003] = 14'b0000000_0000000;
		Dminus[4004] = 14'b0000000_0000000;
		Dminus[4005] = 14'b0000000_0000000;
		Dminus[4006] = 14'b0000000_0000000;
		Dminus[4007] = 14'b0000000_0000000;
		Dminus[4008] = 14'b0000000_0000000;
		Dminus[4009] = 14'b0000000_0000000;
		Dminus[4010] = 14'b0000000_0000000;
		Dminus[4011] = 14'b0000000_0000000;
		Dminus[4012] = 14'b0000000_0000000;
		Dminus[4013] = 14'b0000000_0000000;
		Dminus[4014] = 14'b0000000_0000000;
		Dminus[4015] = 14'b0000000_0000000;
		Dminus[4016] = 14'b0000000_0000000;
		Dminus[4017] = 14'b0000000_0000000;
		Dminus[4018] = 14'b0000000_0000000;
		Dminus[4019] = 14'b0000000_0000000;
		Dminus[4020] = 14'b0000000_0000000;
		Dminus[4021] = 14'b0000000_0000000;
		Dminus[4022] = 14'b0000000_0000000;
		Dminus[4023] = 14'b0000000_0000000;
		Dminus[4024] = 14'b0000000_0000000;
		Dminus[4025] = 14'b0000000_0000000;
		Dminus[4026] = 14'b0000000_0000000;
		Dminus[4027] = 14'b0000000_0000000;
		Dminus[4028] = 14'b0000000_0000000;
		Dminus[4029] = 14'b0000000_0000000;
		Dminus[4030] = 14'b0000000_0000000;
		Dminus[4031] = 14'b0000000_0000000;
		Dminus[4032] = 14'b0000000_0000000;
		Dminus[4033] = 14'b0000000_0000000;
		Dminus[4034] = 14'b0000000_0000000;
		Dminus[4035] = 14'b0000000_0000000;
		Dminus[4036] = 14'b0000000_0000000;
		Dminus[4037] = 14'b0000000_0000000;
		Dminus[4038] = 14'b0000000_0000000;
		Dminus[4039] = 14'b0000000_0000000;
		Dminus[4040] = 14'b0000000_0000000;
		Dminus[4041] = 14'b0000000_0000000;
		Dminus[4042] = 14'b0000000_0000000;
		Dminus[4043] = 14'b0000000_0000000;
		Dminus[4044] = 14'b0000000_0000000;
		Dminus[4045] = 14'b0000000_0000000;
		Dminus[4046] = 14'b0000000_0000000;
		Dminus[4047] = 14'b0000000_0000000;
		Dminus[4048] = 14'b0000000_0000000;
		Dminus[4049] = 14'b0000000_0000000;
		Dminus[4050] = 14'b0000000_0000000;
		Dminus[4051] = 14'b0000000_0000000;
		Dminus[4052] = 14'b0000000_0000000;
		Dminus[4053] = 14'b0000000_0000000;
		Dminus[4054] = 14'b0000000_0000000;
		Dminus[4055] = 14'b0000000_0000000;
		Dminus[4056] = 14'b0000000_0000000;
		Dminus[4057] = 14'b0000000_0000000;
		Dminus[4058] = 14'b0000000_0000000;
		Dminus[4059] = 14'b0000000_0000000;
		Dminus[4060] = 14'b0000000_0000000;
		Dminus[4061] = 14'b0000000_0000000;
		Dminus[4062] = 14'b0000000_0000000;
		Dminus[4063] = 14'b0000000_0000000;
		Dminus[4064] = 14'b0000000_0000000;
		Dminus[4065] = 14'b0000000_0000000;
		Dminus[4066] = 14'b0000000_0000000;
		Dminus[4067] = 14'b0000000_0000000;
		Dminus[4068] = 14'b0000000_0000000;
		Dminus[4069] = 14'b0000000_0000000;
		Dminus[4070] = 14'b0000000_0000000;
		Dminus[4071] = 14'b0000000_0000000;
		Dminus[4072] = 14'b0000000_0000000;
		Dminus[4073] = 14'b0000000_0000000;
		Dminus[4074] = 14'b0000000_0000000;
		Dminus[4075] = 14'b0000000_0000000;
		Dminus[4076] = 14'b0000000_0000000;
		Dminus[4077] = 14'b0000000_0000000;
		Dminus[4078] = 14'b0000000_0000000;
		Dminus[4079] = 14'b0000000_0000000;
		Dminus[4080] = 14'b0000000_0000000;
		Dminus[4081] = 14'b0000000_0000000;
		Dminus[4082] = 14'b0000000_0000000;
		Dminus[4083] = 14'b0000000_0000000;
		Dminus[4084] = 14'b0000000_0000000;
		Dminus[4085] = 14'b0000000_0000000;
		Dminus[4086] = 14'b0000000_0000000;
		Dminus[4087] = 14'b0000000_0000000;
		Dminus[4088] = 14'b0000000_0000000;
		Dminus[4089] = 14'b0000000_0000000;
		Dminus[4090] = 14'b0000000_0000000;
		Dminus[4091] = 14'b0000000_0000000;
		Dminus[4092] = 14'b0000000_0000000;
		Dminus[4093] = 14'b0000000_0000000;
		Dminus[4094] = 14'b0000000_0000000;
		Dminus[4095] = 14'b0000000_0000000;
		Dminus[4096] = 14'b0000000_0000000;
		Dminus[4097] = 14'b0000000_0000000;
		Dminus[4098] = 14'b0000000_0000000;
		Dminus[4099] = 14'b0000000_0000000;
		Dminus[4100] = 14'b0000000_0000000;
		Dminus[4101] = 14'b0000000_0000000;
		Dminus[4102] = 14'b0000000_0000000;
		Dminus[4103] = 14'b0000000_0000000;
		Dminus[4104] = 14'b0000000_0000000;
		Dminus[4105] = 14'b0000000_0000000;
		Dminus[4106] = 14'b0000000_0000000;
		Dminus[4107] = 14'b0000000_0000000;
		Dminus[4108] = 14'b0000000_0000000;
		Dminus[4109] = 14'b0000000_0000000;
		Dminus[4110] = 14'b0000000_0000000;
		Dminus[4111] = 14'b0000000_0000000;
		Dminus[4112] = 14'b0000000_0000000;
		Dminus[4113] = 14'b0000000_0000000;
		Dminus[4114] = 14'b0000000_0000000;
		Dminus[4115] = 14'b0000000_0000000;
		Dminus[4116] = 14'b0000000_0000000;
		Dminus[4117] = 14'b0000000_0000000;
		Dminus[4118] = 14'b0000000_0000000;
		Dminus[4119] = 14'b0000000_0000000;
		Dminus[4120] = 14'b0000000_0000000;
		Dminus[4121] = 14'b0000000_0000000;
		Dminus[4122] = 14'b0000000_0000000;
		Dminus[4123] = 14'b0000000_0000000;
		Dminus[4124] = 14'b0000000_0000000;
		Dminus[4125] = 14'b0000000_0000000;
		Dminus[4126] = 14'b0000000_0000000;
		Dminus[4127] = 14'b0000000_0000000;
		Dminus[4128] = 14'b0000000_0000000;
		Dminus[4129] = 14'b0000000_0000000;
		Dminus[4130] = 14'b0000000_0000000;
		Dminus[4131] = 14'b0000000_0000000;
		Dminus[4132] = 14'b0000000_0000000;
		Dminus[4133] = 14'b0000000_0000000;
		Dminus[4134] = 14'b0000000_0000000;
		Dminus[4135] = 14'b0000000_0000000;
		Dminus[4136] = 14'b0000000_0000000;
		Dminus[4137] = 14'b0000000_0000000;
		Dminus[4138] = 14'b0000000_0000000;
		Dminus[4139] = 14'b0000000_0000000;
		Dminus[4140] = 14'b0000000_0000000;
		Dminus[4141] = 14'b0000000_0000000;
		Dminus[4142] = 14'b0000000_0000000;
		Dminus[4143] = 14'b0000000_0000000;
		Dminus[4144] = 14'b0000000_0000000;
		Dminus[4145] = 14'b0000000_0000000;
		Dminus[4146] = 14'b0000000_0000000;
		Dminus[4147] = 14'b0000000_0000000;
		Dminus[4148] = 14'b0000000_0000000;
		Dminus[4149] = 14'b0000000_0000000;
		Dminus[4150] = 14'b0000000_0000000;
		Dminus[4151] = 14'b0000000_0000000;
		Dminus[4152] = 14'b0000000_0000000;
		Dminus[4153] = 14'b0000000_0000000;
		Dminus[4154] = 14'b0000000_0000000;
		Dminus[4155] = 14'b0000000_0000000;
		Dminus[4156] = 14'b0000000_0000000;
		Dminus[4157] = 14'b0000000_0000000;
		Dminus[4158] = 14'b0000000_0000000;
		Dminus[4159] = 14'b0000000_0000000;
		Dminus[4160] = 14'b0000000_0000000;
		Dminus[4161] = 14'b0000000_0000000;
		Dminus[4162] = 14'b0000000_0000000;
		Dminus[4163] = 14'b0000000_0000000;
		Dminus[4164] = 14'b0000000_0000000;
		Dminus[4165] = 14'b0000000_0000000;
		Dminus[4166] = 14'b0000000_0000000;
		Dminus[4167] = 14'b0000000_0000000;
		Dminus[4168] = 14'b0000000_0000000;
		Dminus[4169] = 14'b0000000_0000000;
		Dminus[4170] = 14'b0000000_0000000;
		Dminus[4171] = 14'b0000000_0000000;
		Dminus[4172] = 14'b0000000_0000000;
		Dminus[4173] = 14'b0000000_0000000;
		Dminus[4174] = 14'b0000000_0000000;
		Dminus[4175] = 14'b0000000_0000000;
		Dminus[4176] = 14'b0000000_0000000;
		Dminus[4177] = 14'b0000000_0000000;
		Dminus[4178] = 14'b0000000_0000000;
		Dminus[4179] = 14'b0000000_0000000;
		Dminus[4180] = 14'b0000000_0000000;
		Dminus[4181] = 14'b0000000_0000000;
		Dminus[4182] = 14'b0000000_0000000;
		Dminus[4183] = 14'b0000000_0000000;
		Dminus[4184] = 14'b0000000_0000000;
		Dminus[4185] = 14'b0000000_0000000;
		Dminus[4186] = 14'b0000000_0000000;
		Dminus[4187] = 14'b0000000_0000000;
		Dminus[4188] = 14'b0000000_0000000;
		Dminus[4189] = 14'b0000000_0000000;
		Dminus[4190] = 14'b0000000_0000000;
		Dminus[4191] = 14'b0000000_0000000;
		Dminus[4192] = 14'b0000000_0000000;
		Dminus[4193] = 14'b0000000_0000000;
		Dminus[4194] = 14'b0000000_0000000;
		Dminus[4195] = 14'b0000000_0000000;
		Dminus[4196] = 14'b0000000_0000000;
		Dminus[4197] = 14'b0000000_0000000;
		Dminus[4198] = 14'b0000000_0000000;
		Dminus[4199] = 14'b0000000_0000000;
		Dminus[4200] = 14'b0000000_0000000;
		Dminus[4201] = 14'b0000000_0000000;
		Dminus[4202] = 14'b0000000_0000000;
		Dminus[4203] = 14'b0000000_0000000;
		Dminus[4204] = 14'b0000000_0000000;
		Dminus[4205] = 14'b0000000_0000000;
		Dminus[4206] = 14'b0000000_0000000;
		Dminus[4207] = 14'b0000000_0000000;
		Dminus[4208] = 14'b0000000_0000000;
		Dminus[4209] = 14'b0000000_0000000;
		Dminus[4210] = 14'b0000000_0000000;
		Dminus[4211] = 14'b0000000_0000000;
		Dminus[4212] = 14'b0000000_0000000;
		Dminus[4213] = 14'b0000000_0000000;
		Dminus[4214] = 14'b0000000_0000000;
		Dminus[4215] = 14'b0000000_0000000;
		Dminus[4216] = 14'b0000000_0000000;
		Dminus[4217] = 14'b0000000_0000000;
		Dminus[4218] = 14'b0000000_0000000;
		Dminus[4219] = 14'b0000000_0000000;
		Dminus[4220] = 14'b0000000_0000000;
		Dminus[4221] = 14'b0000000_0000000;
		Dminus[4222] = 14'b0000000_0000000;
		Dminus[4223] = 14'b0000000_0000000;
		Dminus[4224] = 14'b0000000_0000000;
		Dminus[4225] = 14'b0000000_0000000;
		Dminus[4226] = 14'b0000000_0000000;
		Dminus[4227] = 14'b0000000_0000000;
		Dminus[4228] = 14'b0000000_0000000;
		Dminus[4229] = 14'b0000000_0000000;
		Dminus[4230] = 14'b0000000_0000000;
		Dminus[4231] = 14'b0000000_0000000;
		Dminus[4232] = 14'b0000000_0000000;
		Dminus[4233] = 14'b0000000_0000000;
		Dminus[4234] = 14'b0000000_0000000;
		Dminus[4235] = 14'b0000000_0000000;
		Dminus[4236] = 14'b0000000_0000000;
		Dminus[4237] = 14'b0000000_0000000;
		Dminus[4238] = 14'b0000000_0000000;
		Dminus[4239] = 14'b0000000_0000000;
		Dminus[4240] = 14'b0000000_0000000;
		Dminus[4241] = 14'b0000000_0000000;
		Dminus[4242] = 14'b0000000_0000000;
		Dminus[4243] = 14'b0000000_0000000;
		Dminus[4244] = 14'b0000000_0000000;
		Dminus[4245] = 14'b0000000_0000000;
		Dminus[4246] = 14'b0000000_0000000;
		Dminus[4247] = 14'b0000000_0000000;
		Dminus[4248] = 14'b0000000_0000000;
		Dminus[4249] = 14'b0000000_0000000;
		Dminus[4250] = 14'b0000000_0000000;
		Dminus[4251] = 14'b0000000_0000000;
		Dminus[4252] = 14'b0000000_0000000;
		Dminus[4253] = 14'b0000000_0000000;
		Dminus[4254] = 14'b0000000_0000000;
		Dminus[4255] = 14'b0000000_0000000;
		Dminus[4256] = 14'b0000000_0000000;
		Dminus[4257] = 14'b0000000_0000000;
		Dminus[4258] = 14'b0000000_0000000;
		Dminus[4259] = 14'b0000000_0000000;
		Dminus[4260] = 14'b0000000_0000000;
		Dminus[4261] = 14'b0000000_0000000;
		Dminus[4262] = 14'b0000000_0000000;
		Dminus[4263] = 14'b0000000_0000000;
		Dminus[4264] = 14'b0000000_0000000;
		Dminus[4265] = 14'b0000000_0000000;
		Dminus[4266] = 14'b0000000_0000000;
		Dminus[4267] = 14'b0000000_0000000;
		Dminus[4268] = 14'b0000000_0000000;
		Dminus[4269] = 14'b0000000_0000000;
		Dminus[4270] = 14'b0000000_0000000;
		Dminus[4271] = 14'b0000000_0000000;
		Dminus[4272] = 14'b0000000_0000000;
		Dminus[4273] = 14'b0000000_0000000;
		Dminus[4274] = 14'b0000000_0000000;
		Dminus[4275] = 14'b0000000_0000000;
		Dminus[4276] = 14'b0000000_0000000;
		Dminus[4277] = 14'b0000000_0000000;
		Dminus[4278] = 14'b0000000_0000000;
		Dminus[4279] = 14'b0000000_0000000;
		Dminus[4280] = 14'b0000000_0000000;
		Dminus[4281] = 14'b0000000_0000000;
		Dminus[4282] = 14'b0000000_0000000;
		Dminus[4283] = 14'b0000000_0000000;
		Dminus[4284] = 14'b0000000_0000000;
		Dminus[4285] = 14'b0000000_0000000;
		Dminus[4286] = 14'b0000000_0000000;
		Dminus[4287] = 14'b0000000_0000000;
		Dminus[4288] = 14'b0000000_0000000;
		Dminus[4289] = 14'b0000000_0000000;
		Dminus[4290] = 14'b0000000_0000000;
		Dminus[4291] = 14'b0000000_0000000;
		Dminus[4292] = 14'b0000000_0000000;
		Dminus[4293] = 14'b0000000_0000000;
		Dminus[4294] = 14'b0000000_0000000;
		Dminus[4295] = 14'b0000000_0000000;
		Dminus[4296] = 14'b0000000_0000000;
		Dminus[4297] = 14'b0000000_0000000;
		Dminus[4298] = 14'b0000000_0000000;
		Dminus[4299] = 14'b0000000_0000000;
		Dminus[4300] = 14'b0000000_0000000;
		Dminus[4301] = 14'b0000000_0000000;
		Dminus[4302] = 14'b0000000_0000000;
		Dminus[4303] = 14'b0000000_0000000;
		Dminus[4304] = 14'b0000000_0000000;
		Dminus[4305] = 14'b0000000_0000000;
		Dminus[4306] = 14'b0000000_0000000;
		Dminus[4307] = 14'b0000000_0000000;
		Dminus[4308] = 14'b0000000_0000000;
		Dminus[4309] = 14'b0000000_0000000;
		Dminus[4310] = 14'b0000000_0000000;
		Dminus[4311] = 14'b0000000_0000000;
		Dminus[4312] = 14'b0000000_0000000;
		Dminus[4313] = 14'b0000000_0000000;
		Dminus[4314] = 14'b0000000_0000000;
		Dminus[4315] = 14'b0000000_0000000;
		Dminus[4316] = 14'b0000000_0000000;
		Dminus[4317] = 14'b0000000_0000000;
		Dminus[4318] = 14'b0000000_0000000;
		Dminus[4319] = 14'b0000000_0000000;
		Dminus[4320] = 14'b0000000_0000000;
		Dminus[4321] = 14'b0000000_0000000;
		Dminus[4322] = 14'b0000000_0000000;
		Dminus[4323] = 14'b0000000_0000000;
		Dminus[4324] = 14'b0000000_0000000;
		Dminus[4325] = 14'b0000000_0000000;
		Dminus[4326] = 14'b0000000_0000000;
		Dminus[4327] = 14'b0000000_0000000;
		Dminus[4328] = 14'b0000000_0000000;
		Dminus[4329] = 14'b0000000_0000000;
		Dminus[4330] = 14'b0000000_0000000;
		Dminus[4331] = 14'b0000000_0000000;
		Dminus[4332] = 14'b0000000_0000000;
		Dminus[4333] = 14'b0000000_0000000;
		Dminus[4334] = 14'b0000000_0000000;
		Dminus[4335] = 14'b0000000_0000000;
		Dminus[4336] = 14'b0000000_0000000;
		Dminus[4337] = 14'b0000000_0000000;
		Dminus[4338] = 14'b0000000_0000000;
		Dminus[4339] = 14'b0000000_0000000;
		Dminus[4340] = 14'b0000000_0000000;
		Dminus[4341] = 14'b0000000_0000000;
		Dminus[4342] = 14'b0000000_0000000;
		Dminus[4343] = 14'b0000000_0000000;
		Dminus[4344] = 14'b0000000_0000000;
		Dminus[4345] = 14'b0000000_0000000;
		Dminus[4346] = 14'b0000000_0000000;
		Dminus[4347] = 14'b0000000_0000000;
		Dminus[4348] = 14'b0000000_0000000;
		Dminus[4349] = 14'b0000000_0000000;
		Dminus[4350] = 14'b0000000_0000000;
		Dminus[4351] = 14'b0000000_0000000;
		Dminus[4352] = 14'b0000000_0000000;
		Dminus[4353] = 14'b0000000_0000000;
		Dminus[4354] = 14'b0000000_0000000;
		Dminus[4355] = 14'b0000000_0000000;
		Dminus[4356] = 14'b0000000_0000000;
		Dminus[4357] = 14'b0000000_0000000;
		Dminus[4358] = 14'b0000000_0000000;
		Dminus[4359] = 14'b0000000_0000000;
		Dminus[4360] = 14'b0000000_0000000;
		Dminus[4361] = 14'b0000000_0000000;
		Dminus[4362] = 14'b0000000_0000000;
		Dminus[4363] = 14'b0000000_0000000;
		Dminus[4364] = 14'b0000000_0000000;
		Dminus[4365] = 14'b0000000_0000000;
		Dminus[4366] = 14'b0000000_0000000;
		Dminus[4367] = 14'b0000000_0000000;
		Dminus[4368] = 14'b0000000_0000000;
		Dminus[4369] = 14'b0000000_0000000;
		Dminus[4370] = 14'b0000000_0000000;
		Dminus[4371] = 14'b0000000_0000000;
		Dminus[4372] = 14'b0000000_0000000;
		Dminus[4373] = 14'b0000000_0000000;
		Dminus[4374] = 14'b0000000_0000000;
		Dminus[4375] = 14'b0000000_0000000;
		Dminus[4376] = 14'b0000000_0000000;
		Dminus[4377] = 14'b0000000_0000000;
		Dminus[4378] = 14'b0000000_0000000;
		Dminus[4379] = 14'b0000000_0000000;
		Dminus[4380] = 14'b0000000_0000000;
		Dminus[4381] = 14'b0000000_0000000;
		Dminus[4382] = 14'b0000000_0000000;
		Dminus[4383] = 14'b0000000_0000000;
		Dminus[4384] = 14'b0000000_0000000;
		Dminus[4385] = 14'b0000000_0000000;
		Dminus[4386] = 14'b0000000_0000000;
		Dminus[4387] = 14'b0000000_0000000;
		Dminus[4388] = 14'b0000000_0000000;
		Dminus[4389] = 14'b0000000_0000000;
		Dminus[4390] = 14'b0000000_0000000;
		Dminus[4391] = 14'b0000000_0000000;
		Dminus[4392] = 14'b0000000_0000000;
		Dminus[4393] = 14'b0000000_0000000;
		Dminus[4394] = 14'b0000000_0000000;
		Dminus[4395] = 14'b0000000_0000000;
		Dminus[4396] = 14'b0000000_0000000;
		Dminus[4397] = 14'b0000000_0000000;
		Dminus[4398] = 14'b0000000_0000000;
		Dminus[4399] = 14'b0000000_0000000;
		Dminus[4400] = 14'b0000000_0000000;
		Dminus[4401] = 14'b0000000_0000000;
		Dminus[4402] = 14'b0000000_0000000;
		Dminus[4403] = 14'b0000000_0000000;
		Dminus[4404] = 14'b0000000_0000000;
		Dminus[4405] = 14'b0000000_0000000;
		Dminus[4406] = 14'b0000000_0000000;
		Dminus[4407] = 14'b0000000_0000000;
		Dminus[4408] = 14'b0000000_0000000;
		Dminus[4409] = 14'b0000000_0000000;
		Dminus[4410] = 14'b0000000_0000000;
		Dminus[4411] = 14'b0000000_0000000;
		Dminus[4412] = 14'b0000000_0000000;
		Dminus[4413] = 14'b0000000_0000000;
		Dminus[4414] = 14'b0000000_0000000;
		Dminus[4415] = 14'b0000000_0000000;
		Dminus[4416] = 14'b0000000_0000000;
		Dminus[4417] = 14'b0000000_0000000;
		Dminus[4418] = 14'b0000000_0000000;
		Dminus[4419] = 14'b0000000_0000000;
		Dminus[4420] = 14'b0000000_0000000;
		Dminus[4421] = 14'b0000000_0000000;
		Dminus[4422] = 14'b0000000_0000000;
		Dminus[4423] = 14'b0000000_0000000;
		Dminus[4424] = 14'b0000000_0000000;
		Dminus[4425] = 14'b0000000_0000000;
		Dminus[4426] = 14'b0000000_0000000;
		Dminus[4427] = 14'b0000000_0000000;
		Dminus[4428] = 14'b0000000_0000000;
		Dminus[4429] = 14'b0000000_0000000;
		Dminus[4430] = 14'b0000000_0000000;
		Dminus[4431] = 14'b0000000_0000000;
		Dminus[4432] = 14'b0000000_0000000;
		Dminus[4433] = 14'b0000000_0000000;
		Dminus[4434] = 14'b0000000_0000000;
		Dminus[4435] = 14'b0000000_0000000;
		Dminus[4436] = 14'b0000000_0000000;
		Dminus[4437] = 14'b0000000_0000000;
		Dminus[4438] = 14'b0000000_0000000;
		Dminus[4439] = 14'b0000000_0000000;
		Dminus[4440] = 14'b0000000_0000000;
		Dminus[4441] = 14'b0000000_0000000;
		Dminus[4442] = 14'b0000000_0000000;
		Dminus[4443] = 14'b0000000_0000000;
		Dminus[4444] = 14'b0000000_0000000;
		Dminus[4445] = 14'b0000000_0000000;
		Dminus[4446] = 14'b0000000_0000000;
		Dminus[4447] = 14'b0000000_0000000;
		Dminus[4448] = 14'b0000000_0000000;
		Dminus[4449] = 14'b0000000_0000000;
		Dminus[4450] = 14'b0000000_0000000;
		Dminus[4451] = 14'b0000000_0000000;
		Dminus[4452] = 14'b0000000_0000000;
		Dminus[4453] = 14'b0000000_0000000;
		Dminus[4454] = 14'b0000000_0000000;
		Dminus[4455] = 14'b0000000_0000000;
		Dminus[4456] = 14'b0000000_0000000;
		Dminus[4457] = 14'b0000000_0000000;
		Dminus[4458] = 14'b0000000_0000000;
		Dminus[4459] = 14'b0000000_0000000;
		Dminus[4460] = 14'b0000000_0000000;
		Dminus[4461] = 14'b0000000_0000000;
		Dminus[4462] = 14'b0000000_0000000;
		Dminus[4463] = 14'b0000000_0000000;
		Dminus[4464] = 14'b0000000_0000000;
		Dminus[4465] = 14'b0000000_0000000;
		Dminus[4466] = 14'b0000000_0000000;
		Dminus[4467] = 14'b0000000_0000000;
		Dminus[4468] = 14'b0000000_0000000;
		Dminus[4469] = 14'b0000000_0000000;
		Dminus[4470] = 14'b0000000_0000000;
		Dminus[4471] = 14'b0000000_0000000;
		Dminus[4472] = 14'b0000000_0000000;
		Dminus[4473] = 14'b0000000_0000000;
		Dminus[4474] = 14'b0000000_0000000;
		Dminus[4475] = 14'b0000000_0000000;
		Dminus[4476] = 14'b0000000_0000000;
		Dminus[4477] = 14'b0000000_0000000;
		Dminus[4478] = 14'b0000000_0000000;
		Dminus[4479] = 14'b0000000_0000000;
		Dminus[4480] = 14'b0000000_0000000;
		Dminus[4481] = 14'b0000000_0000000;
		Dminus[4482] = 14'b0000000_0000000;
		Dminus[4483] = 14'b0000000_0000000;
		Dminus[4484] = 14'b0000000_0000000;
		Dminus[4485] = 14'b0000000_0000000;
		Dminus[4486] = 14'b0000000_0000000;
		Dminus[4487] = 14'b0000000_0000000;
		Dminus[4488] = 14'b0000000_0000000;
		Dminus[4489] = 14'b0000000_0000000;
		Dminus[4490] = 14'b0000000_0000000;
		Dminus[4491] = 14'b0000000_0000000;
		Dminus[4492] = 14'b0000000_0000000;
		Dminus[4493] = 14'b0000000_0000000;
		Dminus[4494] = 14'b0000000_0000000;
		Dminus[4495] = 14'b0000000_0000000;
		Dminus[4496] = 14'b0000000_0000000;
		Dminus[4497] = 14'b0000000_0000000;
		Dminus[4498] = 14'b0000000_0000000;
		Dminus[4499] = 14'b0000000_0000000;
		Dminus[4500] = 14'b0000000_0000000;
		Dminus[4501] = 14'b0000000_0000000;
		Dminus[4502] = 14'b0000000_0000000;
		Dminus[4503] = 14'b0000000_0000000;
		Dminus[4504] = 14'b0000000_0000000;
		Dminus[4505] = 14'b0000000_0000000;
		Dminus[4506] = 14'b0000000_0000000;
		Dminus[4507] = 14'b0000000_0000000;
		Dminus[4508] = 14'b0000000_0000000;
		Dminus[4509] = 14'b0000000_0000000;
		Dminus[4510] = 14'b0000000_0000000;
		Dminus[4511] = 14'b0000000_0000000;
		Dminus[4512] = 14'b0000000_0000000;
		Dminus[4513] = 14'b0000000_0000000;
		Dminus[4514] = 14'b0000000_0000000;
		Dminus[4515] = 14'b0000000_0000000;
		Dminus[4516] = 14'b0000000_0000000;
		Dminus[4517] = 14'b0000000_0000000;
		Dminus[4518] = 14'b0000000_0000000;
		Dminus[4519] = 14'b0000000_0000000;
		Dminus[4520] = 14'b0000000_0000000;
		Dminus[4521] = 14'b0000000_0000000;
		Dminus[4522] = 14'b0000000_0000000;
		Dminus[4523] = 14'b0000000_0000000;
		Dminus[4524] = 14'b0000000_0000000;
		Dminus[4525] = 14'b0000000_0000000;
		Dminus[4526] = 14'b0000000_0000000;
		Dminus[4527] = 14'b0000000_0000000;
		Dminus[4528] = 14'b0000000_0000000;
		Dminus[4529] = 14'b0000000_0000000;
		Dminus[4530] = 14'b0000000_0000000;
		Dminus[4531] = 14'b0000000_0000000;
		Dminus[4532] = 14'b0000000_0000000;
		Dminus[4533] = 14'b0000000_0000000;
		Dminus[4534] = 14'b0000000_0000000;
		Dminus[4535] = 14'b0000000_0000000;
		Dminus[4536] = 14'b0000000_0000000;
		Dminus[4537] = 14'b0000000_0000000;
		Dminus[4538] = 14'b0000000_0000000;
		Dminus[4539] = 14'b0000000_0000000;
		Dminus[4540] = 14'b0000000_0000000;
		Dminus[4541] = 14'b0000000_0000000;
		Dminus[4542] = 14'b0000000_0000000;
		Dminus[4543] = 14'b0000000_0000000;
		Dminus[4544] = 14'b0000000_0000000;
		Dminus[4545] = 14'b0000000_0000000;
		Dminus[4546] = 14'b0000000_0000000;
		Dminus[4547] = 14'b0000000_0000000;
		Dminus[4548] = 14'b0000000_0000000;
		Dminus[4549] = 14'b0000000_0000000;
		Dminus[4550] = 14'b0000000_0000000;
		Dminus[4551] = 14'b0000000_0000000;
		Dminus[4552] = 14'b0000000_0000000;
		Dminus[4553] = 14'b0000000_0000000;
		Dminus[4554] = 14'b0000000_0000000;
		Dminus[4555] = 14'b0000000_0000000;
		Dminus[4556] = 14'b0000000_0000000;
		Dminus[4557] = 14'b0000000_0000000;
		Dminus[4558] = 14'b0000000_0000000;
		Dminus[4559] = 14'b0000000_0000000;
		Dminus[4560] = 14'b0000000_0000000;
		Dminus[4561] = 14'b0000000_0000000;
		Dminus[4562] = 14'b0000000_0000000;
		Dminus[4563] = 14'b0000000_0000000;
		Dminus[4564] = 14'b0000000_0000000;
		Dminus[4565] = 14'b0000000_0000000;
		Dminus[4566] = 14'b0000000_0000000;
		Dminus[4567] = 14'b0000000_0000000;
		Dminus[4568] = 14'b0000000_0000000;
		Dminus[4569] = 14'b0000000_0000000;
		Dminus[4570] = 14'b0000000_0000000;
		Dminus[4571] = 14'b0000000_0000000;
		Dminus[4572] = 14'b0000000_0000000;
		Dminus[4573] = 14'b0000000_0000000;
		Dminus[4574] = 14'b0000000_0000000;
		Dminus[4575] = 14'b0000000_0000000;
		Dminus[4576] = 14'b0000000_0000000;
		Dminus[4577] = 14'b0000000_0000000;
		Dminus[4578] = 14'b0000000_0000000;
		Dminus[4579] = 14'b0000000_0000000;
		Dminus[4580] = 14'b0000000_0000000;
		Dminus[4581] = 14'b0000000_0000000;
		Dminus[4582] = 14'b0000000_0000000;
		Dminus[4583] = 14'b0000000_0000000;
		Dminus[4584] = 14'b0000000_0000000;
		Dminus[4585] = 14'b0000000_0000000;
		Dminus[4586] = 14'b0000000_0000000;
		Dminus[4587] = 14'b0000000_0000000;
		Dminus[4588] = 14'b0000000_0000000;
		Dminus[4589] = 14'b0000000_0000000;
		Dminus[4590] = 14'b0000000_0000000;
		Dminus[4591] = 14'b0000000_0000000;
		Dminus[4592] = 14'b0000000_0000000;
		Dminus[4593] = 14'b0000000_0000000;
		Dminus[4594] = 14'b0000000_0000000;
		Dminus[4595] = 14'b0000000_0000000;
		Dminus[4596] = 14'b0000000_0000000;
		Dminus[4597] = 14'b0000000_0000000;
		Dminus[4598] = 14'b0000000_0000000;
		Dminus[4599] = 14'b0000000_0000000;
		Dminus[4600] = 14'b0000000_0000000;
		Dminus[4601] = 14'b0000000_0000000;
		Dminus[4602] = 14'b0000000_0000000;
		Dminus[4603] = 14'b0000000_0000000;
		Dminus[4604] = 14'b0000000_0000000;
		Dminus[4605] = 14'b0000000_0000000;
		Dminus[4606] = 14'b0000000_0000000;
		Dminus[4607] = 14'b0000000_0000000;
		Dminus[4608] = 14'b0000000_0000000;
		Dminus[4609] = 14'b0000000_0000000;
		Dminus[4610] = 14'b0000000_0000000;
		Dminus[4611] = 14'b0000000_0000000;
		Dminus[4612] = 14'b0000000_0000000;
		Dminus[4613] = 14'b0000000_0000000;
		Dminus[4614] = 14'b0000000_0000000;
		Dminus[4615] = 14'b0000000_0000000;
		Dminus[4616] = 14'b0000000_0000000;
		Dminus[4617] = 14'b0000000_0000000;
		Dminus[4618] = 14'b0000000_0000000;
		Dminus[4619] = 14'b0000000_0000000;
		Dminus[4620] = 14'b0000000_0000000;
		Dminus[4621] = 14'b0000000_0000000;
		Dminus[4622] = 14'b0000000_0000000;
		Dminus[4623] = 14'b0000000_0000000;
		Dminus[4624] = 14'b0000000_0000000;
		Dminus[4625] = 14'b0000000_0000000;
		Dminus[4626] = 14'b0000000_0000000;
		Dminus[4627] = 14'b0000000_0000000;
		Dminus[4628] = 14'b0000000_0000000;
		Dminus[4629] = 14'b0000000_0000000;
		Dminus[4630] = 14'b0000000_0000000;
		Dminus[4631] = 14'b0000000_0000000;
		Dminus[4632] = 14'b0000000_0000000;
		Dminus[4633] = 14'b0000000_0000000;
		Dminus[4634] = 14'b0000000_0000000;
		Dminus[4635] = 14'b0000000_0000000;
		Dminus[4636] = 14'b0000000_0000000;
		Dminus[4637] = 14'b0000000_0000000;
		Dminus[4638] = 14'b0000000_0000000;
		Dminus[4639] = 14'b0000000_0000000;
		Dminus[4640] = 14'b0000000_0000000;
		Dminus[4641] = 14'b0000000_0000000;
		Dminus[4642] = 14'b0000000_0000000;
		Dminus[4643] = 14'b0000000_0000000;
		Dminus[4644] = 14'b0000000_0000000;
		Dminus[4645] = 14'b0000000_0000000;
		Dminus[4646] = 14'b0000000_0000000;
		Dminus[4647] = 14'b0000000_0000000;
		Dminus[4648] = 14'b0000000_0000000;
		Dminus[4649] = 14'b0000000_0000000;
		Dminus[4650] = 14'b0000000_0000000;
		Dminus[4651] = 14'b0000000_0000000;
		Dminus[4652] = 14'b0000000_0000000;
		Dminus[4653] = 14'b0000000_0000000;
		Dminus[4654] = 14'b0000000_0000000;
		Dminus[4655] = 14'b0000000_0000000;
		Dminus[4656] = 14'b0000000_0000000;
		Dminus[4657] = 14'b0000000_0000000;
		Dminus[4658] = 14'b0000000_0000000;
		Dminus[4659] = 14'b0000000_0000000;
		Dminus[4660] = 14'b0000000_0000000;
		Dminus[4661] = 14'b0000000_0000000;
		Dminus[4662] = 14'b0000000_0000000;
		Dminus[4663] = 14'b0000000_0000000;
		Dminus[4664] = 14'b0000000_0000000;
		Dminus[4665] = 14'b0000000_0000000;
		Dminus[4666] = 14'b0000000_0000000;
		Dminus[4667] = 14'b0000000_0000000;
		Dminus[4668] = 14'b0000000_0000000;
		Dminus[4669] = 14'b0000000_0000000;
		Dminus[4670] = 14'b0000000_0000000;
		Dminus[4671] = 14'b0000000_0000000;
		Dminus[4672] = 14'b0000000_0000000;
		Dminus[4673] = 14'b0000000_0000000;
		Dminus[4674] = 14'b0000000_0000000;
		Dminus[4675] = 14'b0000000_0000000;
		Dminus[4676] = 14'b0000000_0000000;
		Dminus[4677] = 14'b0000000_0000000;
		Dminus[4678] = 14'b0000000_0000000;
		Dminus[4679] = 14'b0000000_0000000;
		Dminus[4680] = 14'b0000000_0000000;
		Dminus[4681] = 14'b0000000_0000000;
		Dminus[4682] = 14'b0000000_0000000;
		Dminus[4683] = 14'b0000000_0000000;
		Dminus[4684] = 14'b0000000_0000000;
		Dminus[4685] = 14'b0000000_0000000;
		Dminus[4686] = 14'b0000000_0000000;
		Dminus[4687] = 14'b0000000_0000000;
		Dminus[4688] = 14'b0000000_0000000;
		Dminus[4689] = 14'b0000000_0000000;
		Dminus[4690] = 14'b0000000_0000000;
		Dminus[4691] = 14'b0000000_0000000;
		Dminus[4692] = 14'b0000000_0000000;
		Dminus[4693] = 14'b0000000_0000000;
		Dminus[4694] = 14'b0000000_0000000;
		Dminus[4695] = 14'b0000000_0000000;
		Dminus[4696] = 14'b0000000_0000000;
		Dminus[4697] = 14'b0000000_0000000;
		Dminus[4698] = 14'b0000000_0000000;
		Dminus[4699] = 14'b0000000_0000000;
		Dminus[4700] = 14'b0000000_0000000;
		Dminus[4701] = 14'b0000000_0000000;
		Dminus[4702] = 14'b0000000_0000000;
		Dminus[4703] = 14'b0000000_0000000;
		Dminus[4704] = 14'b0000000_0000000;
		Dminus[4705] = 14'b0000000_0000000;
		Dminus[4706] = 14'b0000000_0000000;
		Dminus[4707] = 14'b0000000_0000000;
		Dminus[4708] = 14'b0000000_0000000;
		Dminus[4709] = 14'b0000000_0000000;
		Dminus[4710] = 14'b0000000_0000000;
		Dminus[4711] = 14'b0000000_0000000;
		Dminus[4712] = 14'b0000000_0000000;
		Dminus[4713] = 14'b0000000_0000000;
		Dminus[4714] = 14'b0000000_0000000;
		Dminus[4715] = 14'b0000000_0000000;
		Dminus[4716] = 14'b0000000_0000000;
		Dminus[4717] = 14'b0000000_0000000;
		Dminus[4718] = 14'b0000000_0000000;
		Dminus[4719] = 14'b0000000_0000000;
		Dminus[4720] = 14'b0000000_0000000;
		Dminus[4721] = 14'b0000000_0000000;
		Dminus[4722] = 14'b0000000_0000000;
		Dminus[4723] = 14'b0000000_0000000;
		Dminus[4724] = 14'b0000000_0000000;
		Dminus[4725] = 14'b0000000_0000000;
		Dminus[4726] = 14'b0000000_0000000;
		Dminus[4727] = 14'b0000000_0000000;
		Dminus[4728] = 14'b0000000_0000000;
		Dminus[4729] = 14'b0000000_0000000;
		Dminus[4730] = 14'b0000000_0000000;
		Dminus[4731] = 14'b0000000_0000000;
		Dminus[4732] = 14'b0000000_0000000;
		Dminus[4733] = 14'b0000000_0000000;
		Dminus[4734] = 14'b0000000_0000000;
		Dminus[4735] = 14'b0000000_0000000;
		Dminus[4736] = 14'b0000000_0000000;
		Dminus[4737] = 14'b0000000_0000000;
		Dminus[4738] = 14'b0000000_0000000;
		Dminus[4739] = 14'b0000000_0000000;
		Dminus[4740] = 14'b0000000_0000000;
		Dminus[4741] = 14'b0000000_0000000;
		Dminus[4742] = 14'b0000000_0000000;
		Dminus[4743] = 14'b0000000_0000000;
		Dminus[4744] = 14'b0000000_0000000;
		Dminus[4745] = 14'b0000000_0000000;
		Dminus[4746] = 14'b0000000_0000000;
		Dminus[4747] = 14'b0000000_0000000;
		Dminus[4748] = 14'b0000000_0000000;
		Dminus[4749] = 14'b0000000_0000000;
		Dminus[4750] = 14'b0000000_0000000;
		Dminus[4751] = 14'b0000000_0000000;
		Dminus[4752] = 14'b0000000_0000000;
		Dminus[4753] = 14'b0000000_0000000;
		Dminus[4754] = 14'b0000000_0000000;
		Dminus[4755] = 14'b0000000_0000000;
		Dminus[4756] = 14'b0000000_0000000;
		Dminus[4757] = 14'b0000000_0000000;
		Dminus[4758] = 14'b0000000_0000000;
		Dminus[4759] = 14'b0000000_0000000;
		Dminus[4760] = 14'b0000000_0000000;
		Dminus[4761] = 14'b0000000_0000000;
		Dminus[4762] = 14'b0000000_0000000;
		Dminus[4763] = 14'b0000000_0000000;
		Dminus[4764] = 14'b0000000_0000000;
		Dminus[4765] = 14'b0000000_0000000;
		Dminus[4766] = 14'b0000000_0000000;
		Dminus[4767] = 14'b0000000_0000000;
		Dminus[4768] = 14'b0000000_0000000;
		Dminus[4769] = 14'b0000000_0000000;
		Dminus[4770] = 14'b0000000_0000000;
		Dminus[4771] = 14'b0000000_0000000;
		Dminus[4772] = 14'b0000000_0000000;
		Dminus[4773] = 14'b0000000_0000000;
		Dminus[4774] = 14'b0000000_0000000;
		Dminus[4775] = 14'b0000000_0000000;
		Dminus[4776] = 14'b0000000_0000000;
		Dminus[4777] = 14'b0000000_0000000;
		Dminus[4778] = 14'b0000000_0000000;
		Dminus[4779] = 14'b0000000_0000000;
		Dminus[4780] = 14'b0000000_0000000;
		Dminus[4781] = 14'b0000000_0000000;
		Dminus[4782] = 14'b0000000_0000000;
		Dminus[4783] = 14'b0000000_0000000;
		Dminus[4784] = 14'b0000000_0000000;
		Dminus[4785] = 14'b0000000_0000000;
		Dminus[4786] = 14'b0000000_0000000;
		Dminus[4787] = 14'b0000000_0000000;
		Dminus[4788] = 14'b0000000_0000000;
		Dminus[4789] = 14'b0000000_0000000;
		Dminus[4790] = 14'b0000000_0000000;
		Dminus[4791] = 14'b0000000_0000000;
		Dminus[4792] = 14'b0000000_0000000;
		Dminus[4793] = 14'b0000000_0000000;
		Dminus[4794] = 14'b0000000_0000000;
		Dminus[4795] = 14'b0000000_0000000;
		Dminus[4796] = 14'b0000000_0000000;
		Dminus[4797] = 14'b0000000_0000000;
		Dminus[4798] = 14'b0000000_0000000;
		Dminus[4799] = 14'b0000000_0000000;
		Dminus[4800] = 14'b0000000_0000000;
		Dminus[4801] = 14'b0000000_0000000;
		Dminus[4802] = 14'b0000000_0000000;
		Dminus[4803] = 14'b0000000_0000000;
		Dminus[4804] = 14'b0000000_0000000;
		Dminus[4805] = 14'b0000000_0000000;
		Dminus[4806] = 14'b0000000_0000000;
		Dminus[4807] = 14'b0000000_0000000;
		Dminus[4808] = 14'b0000000_0000000;
		Dminus[4809] = 14'b0000000_0000000;
		Dminus[4810] = 14'b0000000_0000000;
		Dminus[4811] = 14'b0000000_0000000;
		Dminus[4812] = 14'b0000000_0000000;
		Dminus[4813] = 14'b0000000_0000000;
		Dminus[4814] = 14'b0000000_0000000;
		Dminus[4815] = 14'b0000000_0000000;
		Dminus[4816] = 14'b0000000_0000000;
		Dminus[4817] = 14'b0000000_0000000;
		Dminus[4818] = 14'b0000000_0000000;
		Dminus[4819] = 14'b0000000_0000000;
		Dminus[4820] = 14'b0000000_0000000;
		Dminus[4821] = 14'b0000000_0000000;
		Dminus[4822] = 14'b0000000_0000000;
		Dminus[4823] = 14'b0000000_0000000;
		Dminus[4824] = 14'b0000000_0000000;
		Dminus[4825] = 14'b0000000_0000000;
		Dminus[4826] = 14'b0000000_0000000;
		Dminus[4827] = 14'b0000000_0000000;
		Dminus[4828] = 14'b0000000_0000000;
		Dminus[4829] = 14'b0000000_0000000;
		Dminus[4830] = 14'b0000000_0000000;
		Dminus[4831] = 14'b0000000_0000000;
		Dminus[4832] = 14'b0000000_0000000;
		Dminus[4833] = 14'b0000000_0000000;
		Dminus[4834] = 14'b0000000_0000000;
		Dminus[4835] = 14'b0000000_0000000;
		Dminus[4836] = 14'b0000000_0000000;
		Dminus[4837] = 14'b0000000_0000000;
		Dminus[4838] = 14'b0000000_0000000;
		Dminus[4839] = 14'b0000000_0000000;
		Dminus[4840] = 14'b0000000_0000000;
		Dminus[4841] = 14'b0000000_0000000;
		Dminus[4842] = 14'b0000000_0000000;
		Dminus[4843] = 14'b0000000_0000000;
		Dminus[4844] = 14'b0000000_0000000;
		Dminus[4845] = 14'b0000000_0000000;
		Dminus[4846] = 14'b0000000_0000000;
		Dminus[4847] = 14'b0000000_0000000;
		Dminus[4848] = 14'b0000000_0000000;
		Dminus[4849] = 14'b0000000_0000000;
		Dminus[4850] = 14'b0000000_0000000;
		Dminus[4851] = 14'b0000000_0000000;
		Dminus[4852] = 14'b0000000_0000000;
		Dminus[4853] = 14'b0000000_0000000;
		Dminus[4854] = 14'b0000000_0000000;
		Dminus[4855] = 14'b0000000_0000000;
		Dminus[4856] = 14'b0000000_0000000;
		Dminus[4857] = 14'b0000000_0000000;
		Dminus[4858] = 14'b0000000_0000000;
		Dminus[4859] = 14'b0000000_0000000;
		Dminus[4860] = 14'b0000000_0000000;
		Dminus[4861] = 14'b0000000_0000000;
		Dminus[4862] = 14'b0000000_0000000;
		Dminus[4863] = 14'b0000000_0000000;
		Dminus[4864] = 14'b0000000_0000000;
		Dminus[4865] = 14'b0000000_0000000;
		Dminus[4866] = 14'b0000000_0000000;
		Dminus[4867] = 14'b0000000_0000000;
		Dminus[4868] = 14'b0000000_0000000;
		Dminus[4869] = 14'b0000000_0000000;
		Dminus[4870] = 14'b0000000_0000000;
		Dminus[4871] = 14'b0000000_0000000;
		Dminus[4872] = 14'b0000000_0000000;
		Dminus[4873] = 14'b0000000_0000000;
		Dminus[4874] = 14'b0000000_0000000;
		Dminus[4875] = 14'b0000000_0000000;
		Dminus[4876] = 14'b0000000_0000000;
		Dminus[4877] = 14'b0000000_0000000;
		Dminus[4878] = 14'b0000000_0000000;
		Dminus[4879] = 14'b0000000_0000000;
		Dminus[4880] = 14'b0000000_0000000;
		Dminus[4881] = 14'b0000000_0000000;
		Dminus[4882] = 14'b0000000_0000000;
		Dminus[4883] = 14'b0000000_0000000;
		Dminus[4884] = 14'b0000000_0000000;
		Dminus[4885] = 14'b0000000_0000000;
		Dminus[4886] = 14'b0000000_0000000;
		Dminus[4887] = 14'b0000000_0000000;
		Dminus[4888] = 14'b0000000_0000000;
		Dminus[4889] = 14'b0000000_0000000;
		Dminus[4890] = 14'b0000000_0000000;
		Dminus[4891] = 14'b0000000_0000000;
		Dminus[4892] = 14'b0000000_0000000;
		Dminus[4893] = 14'b0000000_0000000;
		Dminus[4894] = 14'b0000000_0000000;
		Dminus[4895] = 14'b0000000_0000000;
		Dminus[4896] = 14'b0000000_0000000;
		Dminus[4897] = 14'b0000000_0000000;
		Dminus[4898] = 14'b0000000_0000000;
		Dminus[4899] = 14'b0000000_0000000;
		Dminus[4900] = 14'b0000000_0000000;
		Dminus[4901] = 14'b0000000_0000000;
		Dminus[4902] = 14'b0000000_0000000;
		Dminus[4903] = 14'b0000000_0000000;
		Dminus[4904] = 14'b0000000_0000000;
		Dminus[4905] = 14'b0000000_0000000;
		Dminus[4906] = 14'b0000000_0000000;
		Dminus[4907] = 14'b0000000_0000000;
		Dminus[4908] = 14'b0000000_0000000;
		Dminus[4909] = 14'b0000000_0000000;
		Dminus[4910] = 14'b0000000_0000000;
		Dminus[4911] = 14'b0000000_0000000;
		Dminus[4912] = 14'b0000000_0000000;
		Dminus[4913] = 14'b0000000_0000000;
		Dminus[4914] = 14'b0000000_0000000;
		Dminus[4915] = 14'b0000000_0000000;
		Dminus[4916] = 14'b0000000_0000000;
		Dminus[4917] = 14'b0000000_0000000;
		Dminus[4918] = 14'b0000000_0000000;
		Dminus[4919] = 14'b0000000_0000000;
		Dminus[4920] = 14'b0000000_0000000;
		Dminus[4921] = 14'b0000000_0000000;
		Dminus[4922] = 14'b0000000_0000000;
		Dminus[4923] = 14'b0000000_0000000;
		Dminus[4924] = 14'b0000000_0000000;
		Dminus[4925] = 14'b0000000_0000000;
		Dminus[4926] = 14'b0000000_0000000;
		Dminus[4927] = 14'b0000000_0000000;
		Dminus[4928] = 14'b0000000_0000000;
		Dminus[4929] = 14'b0000000_0000000;
		Dminus[4930] = 14'b0000000_0000000;
		Dminus[4931] = 14'b0000000_0000000;
		Dminus[4932] = 14'b0000000_0000000;
		Dminus[4933] = 14'b0000000_0000000;
		Dminus[4934] = 14'b0000000_0000000;
		Dminus[4935] = 14'b0000000_0000000;
		Dminus[4936] = 14'b0000000_0000000;
		Dminus[4937] = 14'b0000000_0000000;
		Dminus[4938] = 14'b0000000_0000000;
		Dminus[4939] = 14'b0000000_0000000;
		Dminus[4940] = 14'b0000000_0000000;
		Dminus[4941] = 14'b0000000_0000000;
		Dminus[4942] = 14'b0000000_0000000;
		Dminus[4943] = 14'b0000000_0000000;
		Dminus[4944] = 14'b0000000_0000000;
		Dminus[4945] = 14'b0000000_0000000;
		Dminus[4946] = 14'b0000000_0000000;
		Dminus[4947] = 14'b0000000_0000000;
		Dminus[4948] = 14'b0000000_0000000;
		Dminus[4949] = 14'b0000000_0000000;
		Dminus[4950] = 14'b0000000_0000000;
		Dminus[4951] = 14'b0000000_0000000;
		Dminus[4952] = 14'b0000000_0000000;
		Dminus[4953] = 14'b0000000_0000000;
		Dminus[4954] = 14'b0000000_0000000;
		Dminus[4955] = 14'b0000000_0000000;
		Dminus[4956] = 14'b0000000_0000000;
		Dminus[4957] = 14'b0000000_0000000;
		Dminus[4958] = 14'b0000000_0000000;
		Dminus[4959] = 14'b0000000_0000000;
		Dminus[4960] = 14'b0000000_0000000;
		Dminus[4961] = 14'b0000000_0000000;
		Dminus[4962] = 14'b0000000_0000000;
		Dminus[4963] = 14'b0000000_0000000;
		Dminus[4964] = 14'b0000000_0000000;
		Dminus[4965] = 14'b0000000_0000000;
		Dminus[4966] = 14'b0000000_0000000;
		Dminus[4967] = 14'b0000000_0000000;
		Dminus[4968] = 14'b0000000_0000000;
		Dminus[4969] = 14'b0000000_0000000;
		Dminus[4970] = 14'b0000000_0000000;
		Dminus[4971] = 14'b0000000_0000000;
		Dminus[4972] = 14'b0000000_0000000;
		Dminus[4973] = 14'b0000000_0000000;
		Dminus[4974] = 14'b0000000_0000000;
		Dminus[4975] = 14'b0000000_0000000;
		Dminus[4976] = 14'b0000000_0000000;
		Dminus[4977] = 14'b0000000_0000000;
		Dminus[4978] = 14'b0000000_0000000;
		Dminus[4979] = 14'b0000000_0000000;
		Dminus[4980] = 14'b0000000_0000000;
		Dminus[4981] = 14'b0000000_0000000;
		Dminus[4982] = 14'b0000000_0000000;
		Dminus[4983] = 14'b0000000_0000000;
		Dminus[4984] = 14'b0000000_0000000;
		Dminus[4985] = 14'b0000000_0000000;
		Dminus[4986] = 14'b0000000_0000000;
		Dminus[4987] = 14'b0000000_0000000;
		Dminus[4988] = 14'b0000000_0000000;
		Dminus[4989] = 14'b0000000_0000000;
		Dminus[4990] = 14'b0000000_0000000;
		Dminus[4991] = 14'b0000000_0000000;
		Dminus[4992] = 14'b0000000_0000000;
		Dminus[4993] = 14'b0000000_0000000;
		Dminus[4994] = 14'b0000000_0000000;
		Dminus[4995] = 14'b0000000_0000000;
		Dminus[4996] = 14'b0000000_0000000;
		Dminus[4997] = 14'b0000000_0000000;
		Dminus[4998] = 14'b0000000_0000000;
		Dminus[4999] = 14'b0000000_0000000;
		Dminus[5000] = 14'b0000000_0000000;
		Dminus[5001] = 14'b0000000_0000000;
		Dminus[5002] = 14'b0000000_0000000;
		Dminus[5003] = 14'b0000000_0000000;
		Dminus[5004] = 14'b0000000_0000000;
		Dminus[5005] = 14'b0000000_0000000;
		Dminus[5006] = 14'b0000000_0000000;
		Dminus[5007] = 14'b0000000_0000000;
		Dminus[5008] = 14'b0000000_0000000;
		Dminus[5009] = 14'b0000000_0000000;
		Dminus[5010] = 14'b0000000_0000000;
		Dminus[5011] = 14'b0000000_0000000;
		Dminus[5012] = 14'b0000000_0000000;
		Dminus[5013] = 14'b0000000_0000000;
		Dminus[5014] = 14'b0000000_0000000;
		Dminus[5015] = 14'b0000000_0000000;
		Dminus[5016] = 14'b0000000_0000000;
		Dminus[5017] = 14'b0000000_0000000;
		Dminus[5018] = 14'b0000000_0000000;
		Dminus[5019] = 14'b0000000_0000000;
		Dminus[5020] = 14'b0000000_0000000;
		Dminus[5021] = 14'b0000000_0000000;
		Dminus[5022] = 14'b0000000_0000000;
		Dminus[5023] = 14'b0000000_0000000;
		Dminus[5024] = 14'b0000000_0000000;
		Dminus[5025] = 14'b0000000_0000000;
		Dminus[5026] = 14'b0000000_0000000;
		Dminus[5027] = 14'b0000000_0000000;
		Dminus[5028] = 14'b0000000_0000000;
		Dminus[5029] = 14'b0000000_0000000;
		Dminus[5030] = 14'b0000000_0000000;
		Dminus[5031] = 14'b0000000_0000000;
		Dminus[5032] = 14'b0000000_0000000;
		Dminus[5033] = 14'b0000000_0000000;
		Dminus[5034] = 14'b0000000_0000000;
		Dminus[5035] = 14'b0000000_0000000;
		Dminus[5036] = 14'b0000000_0000000;
		Dminus[5037] = 14'b0000000_0000000;
		Dminus[5038] = 14'b0000000_0000000;
		Dminus[5039] = 14'b0000000_0000000;
		Dminus[5040] = 14'b0000000_0000000;
		Dminus[5041] = 14'b0000000_0000000;
		Dminus[5042] = 14'b0000000_0000000;
		Dminus[5043] = 14'b0000000_0000000;
		Dminus[5044] = 14'b0000000_0000000;
		Dminus[5045] = 14'b0000000_0000000;
		Dminus[5046] = 14'b0000000_0000000;
		Dminus[5047] = 14'b0000000_0000000;
		Dminus[5048] = 14'b0000000_0000000;
		Dminus[5049] = 14'b0000000_0000000;
		Dminus[5050] = 14'b0000000_0000000;
		Dminus[5051] = 14'b0000000_0000000;
		Dminus[5052] = 14'b0000000_0000000;
		Dminus[5053] = 14'b0000000_0000000;
		Dminus[5054] = 14'b0000000_0000000;
		Dminus[5055] = 14'b0000000_0000000;
		Dminus[5056] = 14'b0000000_0000000;
		Dminus[5057] = 14'b0000000_0000000;
		Dminus[5058] = 14'b0000000_0000000;
		Dminus[5059] = 14'b0000000_0000000;
		Dminus[5060] = 14'b0000000_0000000;
		Dminus[5061] = 14'b0000000_0000000;
		Dminus[5062] = 14'b0000000_0000000;
		Dminus[5063] = 14'b0000000_0000000;
		Dminus[5064] = 14'b0000000_0000000;
		Dminus[5065] = 14'b0000000_0000000;
		Dminus[5066] = 14'b0000000_0000000;
		Dminus[5067] = 14'b0000000_0000000;
		Dminus[5068] = 14'b0000000_0000000;
		Dminus[5069] = 14'b0000000_0000000;
		Dminus[5070] = 14'b0000000_0000000;
		Dminus[5071] = 14'b0000000_0000000;
		Dminus[5072] = 14'b0000000_0000000;
		Dminus[5073] = 14'b0000000_0000000;
		Dminus[5074] = 14'b0000000_0000000;
		Dminus[5075] = 14'b0000000_0000000;
		Dminus[5076] = 14'b0000000_0000000;
		Dminus[5077] = 14'b0000000_0000000;
		Dminus[5078] = 14'b0000000_0000000;
		Dminus[5079] = 14'b0000000_0000000;
		Dminus[5080] = 14'b0000000_0000000;
		Dminus[5081] = 14'b0000000_0000000;
		Dminus[5082] = 14'b0000000_0000000;
		Dminus[5083] = 14'b0000000_0000000;
		Dminus[5084] = 14'b0000000_0000000;
		Dminus[5085] = 14'b0000000_0000000;
		Dminus[5086] = 14'b0000000_0000000;
		Dminus[5087] = 14'b0000000_0000000;
		Dminus[5088] = 14'b0000000_0000000;
		Dminus[5089] = 14'b0000000_0000000;
		Dminus[5090] = 14'b0000000_0000000;
		Dminus[5091] = 14'b0000000_0000000;
		Dminus[5092] = 14'b0000000_0000000;
		Dminus[5093] = 14'b0000000_0000000;
		Dminus[5094] = 14'b0000000_0000000;
		Dminus[5095] = 14'b0000000_0000000;
		Dminus[5096] = 14'b0000000_0000000;
		Dminus[5097] = 14'b0000000_0000000;
		Dminus[5098] = 14'b0000000_0000000;
		Dminus[5099] = 14'b0000000_0000000;
		Dminus[5100] = 14'b0000000_0000000;
		Dminus[5101] = 14'b0000000_0000000;
		Dminus[5102] = 14'b0000000_0000000;
		Dminus[5103] = 14'b0000000_0000000;
		Dminus[5104] = 14'b0000000_0000000;
		Dminus[5105] = 14'b0000000_0000000;
		Dminus[5106] = 14'b0000000_0000000;
		Dminus[5107] = 14'b0000000_0000000;
		Dminus[5108] = 14'b0000000_0000000;
		Dminus[5109] = 14'b0000000_0000000;
		Dminus[5110] = 14'b0000000_0000000;
		Dminus[5111] = 14'b0000000_0000000;
		Dminus[5112] = 14'b0000000_0000000;
		Dminus[5113] = 14'b0000000_0000000;
		Dminus[5114] = 14'b0000000_0000000;
		Dminus[5115] = 14'b0000000_0000000;
		Dminus[5116] = 14'b0000000_0000000;
		Dminus[5117] = 14'b0000000_0000000;
		Dminus[5118] = 14'b0000000_0000000;
		Dminus[5119] = 14'b0000000_0000000;
		Dminus[5120] = 14'b0000000_0000000;
		Dminus[5121] = 14'b0000000_0000000;
		Dminus[5122] = 14'b0000000_0000000;
		Dminus[5123] = 14'b0000000_0000000;
		Dminus[5124] = 14'b0000000_0000000;
		Dminus[5125] = 14'b0000000_0000000;
		Dminus[5126] = 14'b0000000_0000000;
		Dminus[5127] = 14'b0000000_0000000;
		Dminus[5128] = 14'b0000000_0000000;
		Dminus[5129] = 14'b0000000_0000000;
		Dminus[5130] = 14'b0000000_0000000;
		Dminus[5131] = 14'b0000000_0000000;
		Dminus[5132] = 14'b0000000_0000000;
		Dminus[5133] = 14'b0000000_0000000;
		Dminus[5134] = 14'b0000000_0000000;
		Dminus[5135] = 14'b0000000_0000000;
		Dminus[5136] = 14'b0000000_0000000;
		Dminus[5137] = 14'b0000000_0000000;
		Dminus[5138] = 14'b0000000_0000000;
		Dminus[5139] = 14'b0000000_0000000;
		Dminus[5140] = 14'b0000000_0000000;
		Dminus[5141] = 14'b0000000_0000000;
		Dminus[5142] = 14'b0000000_0000000;
		Dminus[5143] = 14'b0000000_0000000;
		Dminus[5144] = 14'b0000000_0000000;
		Dminus[5145] = 14'b0000000_0000000;
		Dminus[5146] = 14'b0000000_0000000;
		Dminus[5147] = 14'b0000000_0000000;
		Dminus[5148] = 14'b0000000_0000000;
		Dminus[5149] = 14'b0000000_0000000;
		Dminus[5150] = 14'b0000000_0000000;
		Dminus[5151] = 14'b0000000_0000000;
		Dminus[5152] = 14'b0000000_0000000;
		Dminus[5153] = 14'b0000000_0000000;
		Dminus[5154] = 14'b0000000_0000000;
		Dminus[5155] = 14'b0000000_0000000;
		Dminus[5156] = 14'b0000000_0000000;
		Dminus[5157] = 14'b0000000_0000000;
		Dminus[5158] = 14'b0000000_0000000;
		Dminus[5159] = 14'b0000000_0000000;
		Dminus[5160] = 14'b0000000_0000000;
		Dminus[5161] = 14'b0000000_0000000;
		Dminus[5162] = 14'b0000000_0000000;
		Dminus[5163] = 14'b0000000_0000000;
		Dminus[5164] = 14'b0000000_0000000;
		Dminus[5165] = 14'b0000000_0000000;
		Dminus[5166] = 14'b0000000_0000000;
		Dminus[5167] = 14'b0000000_0000000;
		Dminus[5168] = 14'b0000000_0000000;
		Dminus[5169] = 14'b0000000_0000000;
		Dminus[5170] = 14'b0000000_0000000;
		Dminus[5171] = 14'b0000000_0000000;
		Dminus[5172] = 14'b0000000_0000000;
		Dminus[5173] = 14'b0000000_0000000;
		Dminus[5174] = 14'b0000000_0000000;
		Dminus[5175] = 14'b0000000_0000000;
		Dminus[5176] = 14'b0000000_0000000;
		Dminus[5177] = 14'b0000000_0000000;
		Dminus[5178] = 14'b0000000_0000000;
		Dminus[5179] = 14'b0000000_0000000;
		Dminus[5180] = 14'b0000000_0000000;
		Dminus[5181] = 14'b0000000_0000000;
		Dminus[5182] = 14'b0000000_0000000;
		Dminus[5183] = 14'b0000000_0000000;
		Dminus[5184] = 14'b0000000_0000000;
		Dminus[5185] = 14'b0000000_0000000;
		Dminus[5186] = 14'b0000000_0000000;
		Dminus[5187] = 14'b0000000_0000000;
		Dminus[5188] = 14'b0000000_0000000;
		Dminus[5189] = 14'b0000000_0000000;
		Dminus[5190] = 14'b0000000_0000000;
		Dminus[5191] = 14'b0000000_0000000;
		Dminus[5192] = 14'b0000000_0000000;
		Dminus[5193] = 14'b0000000_0000000;
		Dminus[5194] = 14'b0000000_0000000;
		Dminus[5195] = 14'b0000000_0000000;
		Dminus[5196] = 14'b0000000_0000000;
		Dminus[5197] = 14'b0000000_0000000;
		Dminus[5198] = 14'b0000000_0000000;
		Dminus[5199] = 14'b0000000_0000000;
		Dminus[5200] = 14'b0000000_0000000;
		Dminus[5201] = 14'b0000000_0000000;
		Dminus[5202] = 14'b0000000_0000000;
		Dminus[5203] = 14'b0000000_0000000;
		Dminus[5204] = 14'b0000000_0000000;
		Dminus[5205] = 14'b0000000_0000000;
		Dminus[5206] = 14'b0000000_0000000;
		Dminus[5207] = 14'b0000000_0000000;
		Dminus[5208] = 14'b0000000_0000000;
		Dminus[5209] = 14'b0000000_0000000;
		Dminus[5210] = 14'b0000000_0000000;
		Dminus[5211] = 14'b0000000_0000000;
		Dminus[5212] = 14'b0000000_0000000;
		Dminus[5213] = 14'b0000000_0000000;
		Dminus[5214] = 14'b0000000_0000000;
		Dminus[5215] = 14'b0000000_0000000;
		Dminus[5216] = 14'b0000000_0000000;
		Dminus[5217] = 14'b0000000_0000000;
		Dminus[5218] = 14'b0000000_0000000;
		Dminus[5219] = 14'b0000000_0000000;
		Dminus[5220] = 14'b0000000_0000000;
		Dminus[5221] = 14'b0000000_0000000;
		Dminus[5222] = 14'b0000000_0000000;
		Dminus[5223] = 14'b0000000_0000000;
		Dminus[5224] = 14'b0000000_0000000;
		Dminus[5225] = 14'b0000000_0000000;
		Dminus[5226] = 14'b0000000_0000000;
		Dminus[5227] = 14'b0000000_0000000;
		Dminus[5228] = 14'b0000000_0000000;
		Dminus[5229] = 14'b0000000_0000000;
		Dminus[5230] = 14'b0000000_0000000;
		Dminus[5231] = 14'b0000000_0000000;
		Dminus[5232] = 14'b0000000_0000000;
		Dminus[5233] = 14'b0000000_0000000;
		Dminus[5234] = 14'b0000000_0000000;
		Dminus[5235] = 14'b0000000_0000000;
		Dminus[5236] = 14'b0000000_0000000;
		Dminus[5237] = 14'b0000000_0000000;
		Dminus[5238] = 14'b0000000_0000000;
		Dminus[5239] = 14'b0000000_0000000;
		Dminus[5240] = 14'b0000000_0000000;
		Dminus[5241] = 14'b0000000_0000000;
		Dminus[5242] = 14'b0000000_0000000;
		Dminus[5243] = 14'b0000000_0000000;
		Dminus[5244] = 14'b0000000_0000000;
		Dminus[5245] = 14'b0000000_0000000;
		Dminus[5246] = 14'b0000000_0000000;
		Dminus[5247] = 14'b0000000_0000000;
		Dminus[5248] = 14'b0000000_0000000;
		Dminus[5249] = 14'b0000000_0000000;
		Dminus[5250] = 14'b0000000_0000000;
		Dminus[5251] = 14'b0000000_0000000;
		Dminus[5252] = 14'b0000000_0000000;
		Dminus[5253] = 14'b0000000_0000000;
		Dminus[5254] = 14'b0000000_0000000;
		Dminus[5255] = 14'b0000000_0000000;
		Dminus[5256] = 14'b0000000_0000000;
		Dminus[5257] = 14'b0000000_0000000;
		Dminus[5258] = 14'b0000000_0000000;
		Dminus[5259] = 14'b0000000_0000000;
		Dminus[5260] = 14'b0000000_0000000;
		Dminus[5261] = 14'b0000000_0000000;
		Dminus[5262] = 14'b0000000_0000000;
		Dminus[5263] = 14'b0000000_0000000;
		Dminus[5264] = 14'b0000000_0000000;
		Dminus[5265] = 14'b0000000_0000000;
		Dminus[5266] = 14'b0000000_0000000;
		Dminus[5267] = 14'b0000000_0000000;
		Dminus[5268] = 14'b0000000_0000000;
		Dminus[5269] = 14'b0000000_0000000;
		Dminus[5270] = 14'b0000000_0000000;
		Dminus[5271] = 14'b0000000_0000000;
		Dminus[5272] = 14'b0000000_0000000;
		Dminus[5273] = 14'b0000000_0000000;
		Dminus[5274] = 14'b0000000_0000000;
		Dminus[5275] = 14'b0000000_0000000;
		Dminus[5276] = 14'b0000000_0000000;
		Dminus[5277] = 14'b0000000_0000000;
		Dminus[5278] = 14'b0000000_0000000;
		Dminus[5279] = 14'b0000000_0000000;
		Dminus[5280] = 14'b0000000_0000000;
		Dminus[5281] = 14'b0000000_0000000;
		Dminus[5282] = 14'b0000000_0000000;
		Dminus[5283] = 14'b0000000_0000000;
		Dminus[5284] = 14'b0000000_0000000;
		Dminus[5285] = 14'b0000000_0000000;
		Dminus[5286] = 14'b0000000_0000000;
		Dminus[5287] = 14'b0000000_0000000;
		Dminus[5288] = 14'b0000000_0000000;
		Dminus[5289] = 14'b0000000_0000000;
		Dminus[5290] = 14'b0000000_0000000;
		Dminus[5291] = 14'b0000000_0000000;
		Dminus[5292] = 14'b0000000_0000000;
		Dminus[5293] = 14'b0000000_0000000;
		Dminus[5294] = 14'b0000000_0000000;
		Dminus[5295] = 14'b0000000_0000000;
		Dminus[5296] = 14'b0000000_0000000;
		Dminus[5297] = 14'b0000000_0000000;
		Dminus[5298] = 14'b0000000_0000000;
		Dminus[5299] = 14'b0000000_0000000;
		Dminus[5300] = 14'b0000000_0000000;
		Dminus[5301] = 14'b0000000_0000000;
		Dminus[5302] = 14'b0000000_0000000;
		Dminus[5303] = 14'b0000000_0000000;
		Dminus[5304] = 14'b0000000_0000000;
		Dminus[5305] = 14'b0000000_0000000;
		Dminus[5306] = 14'b0000000_0000000;
		Dminus[5307] = 14'b0000000_0000000;
		Dminus[5308] = 14'b0000000_0000000;
		Dminus[5309] = 14'b0000000_0000000;
		Dminus[5310] = 14'b0000000_0000000;
		Dminus[5311] = 14'b0000000_0000000;
		Dminus[5312] = 14'b0000000_0000000;
		Dminus[5313] = 14'b0000000_0000000;
		Dminus[5314] = 14'b0000000_0000000;
		Dminus[5315] = 14'b0000000_0000000;
		Dminus[5316] = 14'b0000000_0000000;
		Dminus[5317] = 14'b0000000_0000000;
		Dminus[5318] = 14'b0000000_0000000;
		Dminus[5319] = 14'b0000000_0000000;
		Dminus[5320] = 14'b0000000_0000000;
		Dminus[5321] = 14'b0000000_0000000;
		Dminus[5322] = 14'b0000000_0000000;
		Dminus[5323] = 14'b0000000_0000000;
		Dminus[5324] = 14'b0000000_0000000;
		Dminus[5325] = 14'b0000000_0000000;
		Dminus[5326] = 14'b0000000_0000000;
		Dminus[5327] = 14'b0000000_0000000;
		Dminus[5328] = 14'b0000000_0000000;
		Dminus[5329] = 14'b0000000_0000000;
		Dminus[5330] = 14'b0000000_0000000;
		Dminus[5331] = 14'b0000000_0000000;
		Dminus[5332] = 14'b0000000_0000000;
		Dminus[5333] = 14'b0000000_0000000;
		Dminus[5334] = 14'b0000000_0000000;
		Dminus[5335] = 14'b0000000_0000000;
		Dminus[5336] = 14'b0000000_0000000;
		Dminus[5337] = 14'b0000000_0000000;
		Dminus[5338] = 14'b0000000_0000000;
		Dminus[5339] = 14'b0000000_0000000;
		Dminus[5340] = 14'b0000000_0000000;
		Dminus[5341] = 14'b0000000_0000000;
		Dminus[5342] = 14'b0000000_0000000;
		Dminus[5343] = 14'b0000000_0000000;
		Dminus[5344] = 14'b0000000_0000000;
		Dminus[5345] = 14'b0000000_0000000;
		Dminus[5346] = 14'b0000000_0000000;
		Dminus[5347] = 14'b0000000_0000000;
		Dminus[5348] = 14'b0000000_0000000;
		Dminus[5349] = 14'b0000000_0000000;
		Dminus[5350] = 14'b0000000_0000000;
		Dminus[5351] = 14'b0000000_0000000;
		Dminus[5352] = 14'b0000000_0000000;
		Dminus[5353] = 14'b0000000_0000000;
		Dminus[5354] = 14'b0000000_0000000;
		Dminus[5355] = 14'b0000000_0000000;
		Dminus[5356] = 14'b0000000_0000000;
		Dminus[5357] = 14'b0000000_0000000;
		Dminus[5358] = 14'b0000000_0000000;
		Dminus[5359] = 14'b0000000_0000000;
		Dminus[5360] = 14'b0000000_0000000;
		Dminus[5361] = 14'b0000000_0000000;
		Dminus[5362] = 14'b0000000_0000000;
		Dminus[5363] = 14'b0000000_0000000;
		Dminus[5364] = 14'b0000000_0000000;
		Dminus[5365] = 14'b0000000_0000000;
		Dminus[5366] = 14'b0000000_0000000;
		Dminus[5367] = 14'b0000000_0000000;
		Dminus[5368] = 14'b0000000_0000000;
		Dminus[5369] = 14'b0000000_0000000;
		Dminus[5370] = 14'b0000000_0000000;
		Dminus[5371] = 14'b0000000_0000000;
		Dminus[5372] = 14'b0000000_0000000;
		Dminus[5373] = 14'b0000000_0000000;
		Dminus[5374] = 14'b0000000_0000000;
		Dminus[5375] = 14'b0000000_0000000;
		Dminus[5376] = 14'b0000000_0000000;
		Dminus[5377] = 14'b0000000_0000000;
		Dminus[5378] = 14'b0000000_0000000;
		Dminus[5379] = 14'b0000000_0000000;
		Dminus[5380] = 14'b0000000_0000000;
		Dminus[5381] = 14'b0000000_0000000;
		Dminus[5382] = 14'b0000000_0000000;
		Dminus[5383] = 14'b0000000_0000000;
		Dminus[5384] = 14'b0000000_0000000;
		Dminus[5385] = 14'b0000000_0000000;
		Dminus[5386] = 14'b0000000_0000000;
		Dminus[5387] = 14'b0000000_0000000;
		Dminus[5388] = 14'b0000000_0000000;
		Dminus[5389] = 14'b0000000_0000000;
		Dminus[5390] = 14'b0000000_0000000;
		Dminus[5391] = 14'b0000000_0000000;
		Dminus[5392] = 14'b0000000_0000000;
		Dminus[5393] = 14'b0000000_0000000;
		Dminus[5394] = 14'b0000000_0000000;
		Dminus[5395] = 14'b0000000_0000000;
		Dminus[5396] = 14'b0000000_0000000;
		Dminus[5397] = 14'b0000000_0000000;
		Dminus[5398] = 14'b0000000_0000000;
		Dminus[5399] = 14'b0000000_0000000;
		Dminus[5400] = 14'b0000000_0000000;
		Dminus[5401] = 14'b0000000_0000000;
		Dminus[5402] = 14'b0000000_0000000;
		Dminus[5403] = 14'b0000000_0000000;
		Dminus[5404] = 14'b0000000_0000000;
		Dminus[5405] = 14'b0000000_0000000;
		Dminus[5406] = 14'b0000000_0000000;
		Dminus[5407] = 14'b0000000_0000000;
		Dminus[5408] = 14'b0000000_0000000;
		Dminus[5409] = 14'b0000000_0000000;
		Dminus[5410] = 14'b0000000_0000000;
		Dminus[5411] = 14'b0000000_0000000;
		Dminus[5412] = 14'b0000000_0000000;
		Dminus[5413] = 14'b0000000_0000000;
		Dminus[5414] = 14'b0000000_0000000;
		Dminus[5415] = 14'b0000000_0000000;
		Dminus[5416] = 14'b0000000_0000000;
		Dminus[5417] = 14'b0000000_0000000;
		Dminus[5418] = 14'b0000000_0000000;
		Dminus[5419] = 14'b0000000_0000000;
		Dminus[5420] = 14'b0000000_0000000;
		Dminus[5421] = 14'b0000000_0000000;
		Dminus[5422] = 14'b0000000_0000000;
		Dminus[5423] = 14'b0000000_0000000;
		Dminus[5424] = 14'b0000000_0000000;
		Dminus[5425] = 14'b0000000_0000000;
		Dminus[5426] = 14'b0000000_0000000;
		Dminus[5427] = 14'b0000000_0000000;
		Dminus[5428] = 14'b0000000_0000000;
		Dminus[5429] = 14'b0000000_0000000;
		Dminus[5430] = 14'b0000000_0000000;
		Dminus[5431] = 14'b0000000_0000000;
		Dminus[5432] = 14'b0000000_0000000;
		Dminus[5433] = 14'b0000000_0000000;
		Dminus[5434] = 14'b0000000_0000000;
		Dminus[5435] = 14'b0000000_0000000;
		Dminus[5436] = 14'b0000000_0000000;
		Dminus[5437] = 14'b0000000_0000000;
		Dminus[5438] = 14'b0000000_0000000;
		Dminus[5439] = 14'b0000000_0000000;
		Dminus[5440] = 14'b0000000_0000000;
		Dminus[5441] = 14'b0000000_0000000;
		Dminus[5442] = 14'b0000000_0000000;
		Dminus[5443] = 14'b0000000_0000000;
		Dminus[5444] = 14'b0000000_0000000;
		Dminus[5445] = 14'b0000000_0000000;
		Dminus[5446] = 14'b0000000_0000000;
		Dminus[5447] = 14'b0000000_0000000;
		Dminus[5448] = 14'b0000000_0000000;
		Dminus[5449] = 14'b0000000_0000000;
		Dminus[5450] = 14'b0000000_0000000;
		Dminus[5451] = 14'b0000000_0000000;
		Dminus[5452] = 14'b0000000_0000000;
		Dminus[5453] = 14'b0000000_0000000;
		Dminus[5454] = 14'b0000000_0000000;
		Dminus[5455] = 14'b0000000_0000000;
		Dminus[5456] = 14'b0000000_0000000;
		Dminus[5457] = 14'b0000000_0000000;
		Dminus[5458] = 14'b0000000_0000000;
		Dminus[5459] = 14'b0000000_0000000;
		Dminus[5460] = 14'b0000000_0000000;
		Dminus[5461] = 14'b0000000_0000000;
		Dminus[5462] = 14'b0000000_0000000;
		Dminus[5463] = 14'b0000000_0000000;
		Dminus[5464] = 14'b0000000_0000000;
		Dminus[5465] = 14'b0000000_0000000;
		Dminus[5466] = 14'b0000000_0000000;
		Dminus[5467] = 14'b0000000_0000000;
		Dminus[5468] = 14'b0000000_0000000;
		Dminus[5469] = 14'b0000000_0000000;
		Dminus[5470] = 14'b0000000_0000000;
		Dminus[5471] = 14'b0000000_0000000;
		Dminus[5472] = 14'b0000000_0000000;
		Dminus[5473] = 14'b0000000_0000000;
		Dminus[5474] = 14'b0000000_0000000;
		Dminus[5475] = 14'b0000000_0000000;
		Dminus[5476] = 14'b0000000_0000000;
		Dminus[5477] = 14'b0000000_0000000;
		Dminus[5478] = 14'b0000000_0000000;
		Dminus[5479] = 14'b0000000_0000000;
		Dminus[5480] = 14'b0000000_0000000;
		Dminus[5481] = 14'b0000000_0000000;
		Dminus[5482] = 14'b0000000_0000000;
		Dminus[5483] = 14'b0000000_0000000;
		Dminus[5484] = 14'b0000000_0000000;
		Dminus[5485] = 14'b0000000_0000000;
		Dminus[5486] = 14'b0000000_0000000;
		Dminus[5487] = 14'b0000000_0000000;
		Dminus[5488] = 14'b0000000_0000000;
		Dminus[5489] = 14'b0000000_0000000;
		Dminus[5490] = 14'b0000000_0000000;
		Dminus[5491] = 14'b0000000_0000000;
		Dminus[5492] = 14'b0000000_0000000;
		Dminus[5493] = 14'b0000000_0000000;
		Dminus[5494] = 14'b0000000_0000000;
		Dminus[5495] = 14'b0000000_0000000;
		Dminus[5496] = 14'b0000000_0000000;
		Dminus[5497] = 14'b0000000_0000000;
		Dminus[5498] = 14'b0000000_0000000;
		Dminus[5499] = 14'b0000000_0000000;
		Dminus[5500] = 14'b0000000_0000000;
		Dminus[5501] = 14'b0000000_0000000;
		Dminus[5502] = 14'b0000000_0000000;
		Dminus[5503] = 14'b0000000_0000000;
		Dminus[5504] = 14'b0000000_0000000;
		Dminus[5505] = 14'b0000000_0000000;
		Dminus[5506] = 14'b0000000_0000000;
		Dminus[5507] = 14'b0000000_0000000;
		Dminus[5508] = 14'b0000000_0000000;
		Dminus[5509] = 14'b0000000_0000000;
		Dminus[5510] = 14'b0000000_0000000;
		Dminus[5511] = 14'b0000000_0000000;
		Dminus[5512] = 14'b0000000_0000000;
		Dminus[5513] = 14'b0000000_0000000;
		Dminus[5514] = 14'b0000000_0000000;
		Dminus[5515] = 14'b0000000_0000000;
		Dminus[5516] = 14'b0000000_0000000;
		Dminus[5517] = 14'b0000000_0000000;
		Dminus[5518] = 14'b0000000_0000000;
		Dminus[5519] = 14'b0000000_0000000;
		Dminus[5520] = 14'b0000000_0000000;
		Dminus[5521] = 14'b0000000_0000000;
		Dminus[5522] = 14'b0000000_0000000;
		Dminus[5523] = 14'b0000000_0000000;
		Dminus[5524] = 14'b0000000_0000000;
		Dminus[5525] = 14'b0000000_0000000;
		Dminus[5526] = 14'b0000000_0000000;
		Dminus[5527] = 14'b0000000_0000000;
		Dminus[5528] = 14'b0000000_0000000;
		Dminus[5529] = 14'b0000000_0000000;
		Dminus[5530] = 14'b0000000_0000000;
		Dminus[5531] = 14'b0000000_0000000;
		Dminus[5532] = 14'b0000000_0000000;
		Dminus[5533] = 14'b0000000_0000000;
		Dminus[5534] = 14'b0000000_0000000;
		Dminus[5535] = 14'b0000000_0000000;
		Dminus[5536] = 14'b0000000_0000000;
		Dminus[5537] = 14'b0000000_0000000;
		Dminus[5538] = 14'b0000000_0000000;
		Dminus[5539] = 14'b0000000_0000000;
		Dminus[5540] = 14'b0000000_0000000;
		Dminus[5541] = 14'b0000000_0000000;
		Dminus[5542] = 14'b0000000_0000000;
		Dminus[5543] = 14'b0000000_0000000;
		Dminus[5544] = 14'b0000000_0000000;
		Dminus[5545] = 14'b0000000_0000000;
		Dminus[5546] = 14'b0000000_0000000;
		Dminus[5547] = 14'b0000000_0000000;
		Dminus[5548] = 14'b0000000_0000000;
		Dminus[5549] = 14'b0000000_0000000;
		Dminus[5550] = 14'b0000000_0000000;
		Dminus[5551] = 14'b0000000_0000000;
		Dminus[5552] = 14'b0000000_0000000;
		Dminus[5553] = 14'b0000000_0000000;
		Dminus[5554] = 14'b0000000_0000000;
		Dminus[5555] = 14'b0000000_0000000;
		Dminus[5556] = 14'b0000000_0000000;
		Dminus[5557] = 14'b0000000_0000000;
		Dminus[5558] = 14'b0000000_0000000;
		Dminus[5559] = 14'b0000000_0000000;
		Dminus[5560] = 14'b0000000_0000000;
		Dminus[5561] = 14'b0000000_0000000;
		Dminus[5562] = 14'b0000000_0000000;
		Dminus[5563] = 14'b0000000_0000000;
		Dminus[5564] = 14'b0000000_0000000;
		Dminus[5565] = 14'b0000000_0000000;
		Dminus[5566] = 14'b0000000_0000000;
		Dminus[5567] = 14'b0000000_0000000;
		Dminus[5568] = 14'b0000000_0000000;
		Dminus[5569] = 14'b0000000_0000000;
		Dminus[5570] = 14'b0000000_0000000;
		Dminus[5571] = 14'b0000000_0000000;
		Dminus[5572] = 14'b0000000_0000000;
		Dminus[5573] = 14'b0000000_0000000;
		Dminus[5574] = 14'b0000000_0000000;
		Dminus[5575] = 14'b0000000_0000000;
		Dminus[5576] = 14'b0000000_0000000;
		Dminus[5577] = 14'b0000000_0000000;
		Dminus[5578] = 14'b0000000_0000000;
		Dminus[5579] = 14'b0000000_0000000;
		Dminus[5580] = 14'b0000000_0000000;
		Dminus[5581] = 14'b0000000_0000000;
		Dminus[5582] = 14'b0000000_0000000;
		Dminus[5583] = 14'b0000000_0000000;
		Dminus[5584] = 14'b0000000_0000000;
		Dminus[5585] = 14'b0000000_0000000;
		Dminus[5586] = 14'b0000000_0000000;
		Dminus[5587] = 14'b0000000_0000000;
		Dminus[5588] = 14'b0000000_0000000;
		Dminus[5589] = 14'b0000000_0000000;
		Dminus[5590] = 14'b0000000_0000000;
		Dminus[5591] = 14'b0000000_0000000;
		Dminus[5592] = 14'b0000000_0000000;
		Dminus[5593] = 14'b0000000_0000000;
		Dminus[5594] = 14'b0000000_0000000;
		Dminus[5595] = 14'b0000000_0000000;
		Dminus[5596] = 14'b0000000_0000000;
		Dminus[5597] = 14'b0000000_0000000;
		Dminus[5598] = 14'b0000000_0000000;
		Dminus[5599] = 14'b0000000_0000000;
		Dminus[5600] = 14'b0000000_0000000;
		Dminus[5601] = 14'b0000000_0000000;
		Dminus[5602] = 14'b0000000_0000000;
		Dminus[5603] = 14'b0000000_0000000;
		Dminus[5604] = 14'b0000000_0000000;
		Dminus[5605] = 14'b0000000_0000000;
		Dminus[5606] = 14'b0000000_0000000;
		Dminus[5607] = 14'b0000000_0000000;
		Dminus[5608] = 14'b0000000_0000000;
		Dminus[5609] = 14'b0000000_0000000;
		Dminus[5610] = 14'b0000000_0000000;
		Dminus[5611] = 14'b0000000_0000000;
		Dminus[5612] = 14'b0000000_0000000;
		Dminus[5613] = 14'b0000000_0000000;
		Dminus[5614] = 14'b0000000_0000000;
		Dminus[5615] = 14'b0000000_0000000;
		Dminus[5616] = 14'b0000000_0000000;
		Dminus[5617] = 14'b0000000_0000000;
		Dminus[5618] = 14'b0000000_0000000;
		Dminus[5619] = 14'b0000000_0000000;
		Dminus[5620] = 14'b0000000_0000000;
		Dminus[5621] = 14'b0000000_0000000;
		Dminus[5622] = 14'b0000000_0000000;
		Dminus[5623] = 14'b0000000_0000000;
		Dminus[5624] = 14'b0000000_0000000;
		Dminus[5625] = 14'b0000000_0000000;
		Dminus[5626] = 14'b0000000_0000000;
		Dminus[5627] = 14'b0000000_0000000;
		Dminus[5628] = 14'b0000000_0000000;
		Dminus[5629] = 14'b0000000_0000000;
		Dminus[5630] = 14'b0000000_0000000;
		Dminus[5631] = 14'b0000000_0000000;
		Dminus[5632] = 14'b0000000_0000000;
		Dminus[5633] = 14'b0000000_0000000;
		Dminus[5634] = 14'b0000000_0000000;
		Dminus[5635] = 14'b0000000_0000000;
		Dminus[5636] = 14'b0000000_0000000;
		Dminus[5637] = 14'b0000000_0000000;
		Dminus[5638] = 14'b0000000_0000000;
		Dminus[5639] = 14'b0000000_0000000;
		Dminus[5640] = 14'b0000000_0000000;
		Dminus[5641] = 14'b0000000_0000000;
		Dminus[5642] = 14'b0000000_0000000;
		Dminus[5643] = 14'b0000000_0000000;
		Dminus[5644] = 14'b0000000_0000000;
		Dminus[5645] = 14'b0000000_0000000;
		Dminus[5646] = 14'b0000000_0000000;
		Dminus[5647] = 14'b0000000_0000000;
		Dminus[5648] = 14'b0000000_0000000;
		Dminus[5649] = 14'b0000000_0000000;
		Dminus[5650] = 14'b0000000_0000000;
		Dminus[5651] = 14'b0000000_0000000;
		Dminus[5652] = 14'b0000000_0000000;
		Dminus[5653] = 14'b0000000_0000000;
		Dminus[5654] = 14'b0000000_0000000;
		Dminus[5655] = 14'b0000000_0000000;
		Dminus[5656] = 14'b0000000_0000000;
		Dminus[5657] = 14'b0000000_0000000;
		Dminus[5658] = 14'b0000000_0000000;
		Dminus[5659] = 14'b0000000_0000000;
		Dminus[5660] = 14'b0000000_0000000;
		Dminus[5661] = 14'b0000000_0000000;
		Dminus[5662] = 14'b0000000_0000000;
		Dminus[5663] = 14'b0000000_0000000;
		Dminus[5664] = 14'b0000000_0000000;
		Dminus[5665] = 14'b0000000_0000000;
		Dminus[5666] = 14'b0000000_0000000;
		Dminus[5667] = 14'b0000000_0000000;
		Dminus[5668] = 14'b0000000_0000000;
		Dminus[5669] = 14'b0000000_0000000;
		Dminus[5670] = 14'b0000000_0000000;
		Dminus[5671] = 14'b0000000_0000000;
		Dminus[5672] = 14'b0000000_0000000;
		Dminus[5673] = 14'b0000000_0000000;
		Dminus[5674] = 14'b0000000_0000000;
		Dminus[5675] = 14'b0000000_0000000;
		Dminus[5676] = 14'b0000000_0000000;
		Dminus[5677] = 14'b0000000_0000000;
		Dminus[5678] = 14'b0000000_0000000;
		Dminus[5679] = 14'b0000000_0000000;
		Dminus[5680] = 14'b0000000_0000000;
		Dminus[5681] = 14'b0000000_0000000;
		Dminus[5682] = 14'b0000000_0000000;
		Dminus[5683] = 14'b0000000_0000000;
		Dminus[5684] = 14'b0000000_0000000;
		Dminus[5685] = 14'b0000000_0000000;
		Dminus[5686] = 14'b0000000_0000000;
		Dminus[5687] = 14'b0000000_0000000;
		Dminus[5688] = 14'b0000000_0000000;
		Dminus[5689] = 14'b0000000_0000000;
		Dminus[5690] = 14'b0000000_0000000;
		Dminus[5691] = 14'b0000000_0000000;
		Dminus[5692] = 14'b0000000_0000000;
		Dminus[5693] = 14'b0000000_0000000;
		Dminus[5694] = 14'b0000000_0000000;
		Dminus[5695] = 14'b0000000_0000000;
		Dminus[5696] = 14'b0000000_0000000;
		Dminus[5697] = 14'b0000000_0000000;
		Dminus[5698] = 14'b0000000_0000000;
		Dminus[5699] = 14'b0000000_0000000;
		Dminus[5700] = 14'b0000000_0000000;
		Dminus[5701] = 14'b0000000_0000000;
		Dminus[5702] = 14'b0000000_0000000;
		Dminus[5703] = 14'b0000000_0000000;
		Dminus[5704] = 14'b0000000_0000000;
		Dminus[5705] = 14'b0000000_0000000;
		Dminus[5706] = 14'b0000000_0000000;
		Dminus[5707] = 14'b0000000_0000000;
		Dminus[5708] = 14'b0000000_0000000;
		Dminus[5709] = 14'b0000000_0000000;
		Dminus[5710] = 14'b0000000_0000000;
		Dminus[5711] = 14'b0000000_0000000;
		Dminus[5712] = 14'b0000000_0000000;
		Dminus[5713] = 14'b0000000_0000000;
		Dminus[5714] = 14'b0000000_0000000;
		Dminus[5715] = 14'b0000000_0000000;
		Dminus[5716] = 14'b0000000_0000000;
		Dminus[5717] = 14'b0000000_0000000;
		Dminus[5718] = 14'b0000000_0000000;
		Dminus[5719] = 14'b0000000_0000000;
		Dminus[5720] = 14'b0000000_0000000;
		Dminus[5721] = 14'b0000000_0000000;
		Dminus[5722] = 14'b0000000_0000000;
		Dminus[5723] = 14'b0000000_0000000;
		Dminus[5724] = 14'b0000000_0000000;
		Dminus[5725] = 14'b0000000_0000000;
		Dminus[5726] = 14'b0000000_0000000;
		Dminus[5727] = 14'b0000000_0000000;
		Dminus[5728] = 14'b0000000_0000000;
		Dminus[5729] = 14'b0000000_0000000;
		Dminus[5730] = 14'b0000000_0000000;
		Dminus[5731] = 14'b0000000_0000000;
		Dminus[5732] = 14'b0000000_0000000;
		Dminus[5733] = 14'b0000000_0000000;
		Dminus[5734] = 14'b0000000_0000000;
		Dminus[5735] = 14'b0000000_0000000;
		Dminus[5736] = 14'b0000000_0000000;
		Dminus[5737] = 14'b0000000_0000000;
		Dminus[5738] = 14'b0000000_0000000;
		Dminus[5739] = 14'b0000000_0000000;
		Dminus[5740] = 14'b0000000_0000000;
		Dminus[5741] = 14'b0000000_0000000;
		Dminus[5742] = 14'b0000000_0000000;
		Dminus[5743] = 14'b0000000_0000000;
		Dminus[5744] = 14'b0000000_0000000;
		Dminus[5745] = 14'b0000000_0000000;
		Dminus[5746] = 14'b0000000_0000000;
		Dminus[5747] = 14'b0000000_0000000;
		Dminus[5748] = 14'b0000000_0000000;
		Dminus[5749] = 14'b0000000_0000000;
		Dminus[5750] = 14'b0000000_0000000;
		Dminus[5751] = 14'b0000000_0000000;
		Dminus[5752] = 14'b0000000_0000000;
		Dminus[5753] = 14'b0000000_0000000;
		Dminus[5754] = 14'b0000000_0000000;
		Dminus[5755] = 14'b0000000_0000000;
		Dminus[5756] = 14'b0000000_0000000;
		Dminus[5757] = 14'b0000000_0000000;
		Dminus[5758] = 14'b0000000_0000000;
		Dminus[5759] = 14'b0000000_0000000;
		Dminus[5760] = 14'b0000000_0000000;
		Dminus[5761] = 14'b0000000_0000000;
		Dminus[5762] = 14'b0000000_0000000;
		Dminus[5763] = 14'b0000000_0000000;
		Dminus[5764] = 14'b0000000_0000000;
		Dminus[5765] = 14'b0000000_0000000;
		Dminus[5766] = 14'b0000000_0000000;
		Dminus[5767] = 14'b0000000_0000000;
		Dminus[5768] = 14'b0000000_0000000;
		Dminus[5769] = 14'b0000000_0000000;
		Dminus[5770] = 14'b0000000_0000000;
		Dminus[5771] = 14'b0000000_0000000;
		Dminus[5772] = 14'b0000000_0000000;
		Dminus[5773] = 14'b0000000_0000000;
		Dminus[5774] = 14'b0000000_0000000;
		Dminus[5775] = 14'b0000000_0000000;
		Dminus[5776] = 14'b0000000_0000000;
		Dminus[5777] = 14'b0000000_0000000;
		Dminus[5778] = 14'b0000000_0000000;
		Dminus[5779] = 14'b0000000_0000000;
		Dminus[5780] = 14'b0000000_0000000;
		Dminus[5781] = 14'b0000000_0000000;
		Dminus[5782] = 14'b0000000_0000000;
		Dminus[5783] = 14'b0000000_0000000;
		Dminus[5784] = 14'b0000000_0000000;
		Dminus[5785] = 14'b0000000_0000000;
		Dminus[5786] = 14'b0000000_0000000;
		Dminus[5787] = 14'b0000000_0000000;
		Dminus[5788] = 14'b0000000_0000000;
		Dminus[5789] = 14'b0000000_0000000;
		Dminus[5790] = 14'b0000000_0000000;
		Dminus[5791] = 14'b0000000_0000000;
		Dminus[5792] = 14'b0000000_0000000;
		Dminus[5793] = 14'b0000000_0000000;
		Dminus[5794] = 14'b0000000_0000000;
		Dminus[5795] = 14'b0000000_0000000;
		Dminus[5796] = 14'b0000000_0000000;
		Dminus[5797] = 14'b0000000_0000000;
		Dminus[5798] = 14'b0000000_0000000;
		Dminus[5799] = 14'b0000000_0000000;
		Dminus[5800] = 14'b0000000_0000000;
		Dminus[5801] = 14'b0000000_0000000;
		Dminus[5802] = 14'b0000000_0000000;
		Dminus[5803] = 14'b0000000_0000000;
		Dminus[5804] = 14'b0000000_0000000;
		Dminus[5805] = 14'b0000000_0000000;
		Dminus[5806] = 14'b0000000_0000000;
		Dminus[5807] = 14'b0000000_0000000;
		Dminus[5808] = 14'b0000000_0000000;
		Dminus[5809] = 14'b0000000_0000000;
		Dminus[5810] = 14'b0000000_0000000;
		Dminus[5811] = 14'b0000000_0000000;
		Dminus[5812] = 14'b0000000_0000000;
		Dminus[5813] = 14'b0000000_0000000;
		Dminus[5814] = 14'b0000000_0000000;
		Dminus[5815] = 14'b0000000_0000000;
		Dminus[5816] = 14'b0000000_0000000;
		Dminus[5817] = 14'b0000000_0000000;
		Dminus[5818] = 14'b0000000_0000000;
		Dminus[5819] = 14'b0000000_0000000;
		Dminus[5820] = 14'b0000000_0000000;
		Dminus[5821] = 14'b0000000_0000000;
		Dminus[5822] = 14'b0000000_0000000;
		Dminus[5823] = 14'b0000000_0000000;
		Dminus[5824] = 14'b0000000_0000000;
		Dminus[5825] = 14'b0000000_0000000;
		Dminus[5826] = 14'b0000000_0000000;
		Dminus[5827] = 14'b0000000_0000000;
		Dminus[5828] = 14'b0000000_0000000;
		Dminus[5829] = 14'b0000000_0000000;
		Dminus[5830] = 14'b0000000_0000000;
		Dminus[5831] = 14'b0000000_0000000;
		Dminus[5832] = 14'b0000000_0000000;
		Dminus[5833] = 14'b0000000_0000000;
		Dminus[5834] = 14'b0000000_0000000;
		Dminus[5835] = 14'b0000000_0000000;
		Dminus[5836] = 14'b0000000_0000000;
		Dminus[5837] = 14'b0000000_0000000;
		Dminus[5838] = 14'b0000000_0000000;
		Dminus[5839] = 14'b0000000_0000000;
		Dminus[5840] = 14'b0000000_0000000;
		Dminus[5841] = 14'b0000000_0000000;
		Dminus[5842] = 14'b0000000_0000000;
		Dminus[5843] = 14'b0000000_0000000;
		Dminus[5844] = 14'b0000000_0000000;
		Dminus[5845] = 14'b0000000_0000000;
		Dminus[5846] = 14'b0000000_0000000;
		Dminus[5847] = 14'b0000000_0000000;
		Dminus[5848] = 14'b0000000_0000000;
		Dminus[5849] = 14'b0000000_0000000;
		Dminus[5850] = 14'b0000000_0000000;
		Dminus[5851] = 14'b0000000_0000000;
		Dminus[5852] = 14'b0000000_0000000;
		Dminus[5853] = 14'b0000000_0000000;
		Dminus[5854] = 14'b0000000_0000000;
		Dminus[5855] = 14'b0000000_0000000;
		Dminus[5856] = 14'b0000000_0000000;
		Dminus[5857] = 14'b0000000_0000000;
		Dminus[5858] = 14'b0000000_0000000;
		Dminus[5859] = 14'b0000000_0000000;
		Dminus[5860] = 14'b0000000_0000000;
		Dminus[5861] = 14'b0000000_0000000;
		Dminus[5862] = 14'b0000000_0000000;
		Dminus[5863] = 14'b0000000_0000000;
		Dminus[5864] = 14'b0000000_0000000;
		Dminus[5865] = 14'b0000000_0000000;
		Dminus[5866] = 14'b0000000_0000000;
		Dminus[5867] = 14'b0000000_0000000;
		Dminus[5868] = 14'b0000000_0000000;
		Dminus[5869] = 14'b0000000_0000000;
		Dminus[5870] = 14'b0000000_0000000;
		Dminus[5871] = 14'b0000000_0000000;
		Dminus[5872] = 14'b0000000_0000000;
		Dminus[5873] = 14'b0000000_0000000;
		Dminus[5874] = 14'b0000000_0000000;
		Dminus[5875] = 14'b0000000_0000000;
		Dminus[5876] = 14'b0000000_0000000;
		Dminus[5877] = 14'b0000000_0000000;
		Dminus[5878] = 14'b0000000_0000000;
		Dminus[5879] = 14'b0000000_0000000;
		Dminus[5880] = 14'b0000000_0000000;
		Dminus[5881] = 14'b0000000_0000000;
		Dminus[5882] = 14'b0000000_0000000;
		Dminus[5883] = 14'b0000000_0000000;
		Dminus[5884] = 14'b0000000_0000000;
		Dminus[5885] = 14'b0000000_0000000;
		Dminus[5886] = 14'b0000000_0000000;
		Dminus[5887] = 14'b0000000_0000000;
		Dminus[5888] = 14'b0000000_0000000;
		Dminus[5889] = 14'b0000000_0000000;
		Dminus[5890] = 14'b0000000_0000000;
		Dminus[5891] = 14'b0000000_0000000;
		Dminus[5892] = 14'b0000000_0000000;
		Dminus[5893] = 14'b0000000_0000000;
		Dminus[5894] = 14'b0000000_0000000;
		Dminus[5895] = 14'b0000000_0000000;
		Dminus[5896] = 14'b0000000_0000000;
		Dminus[5897] = 14'b0000000_0000000;
		Dminus[5898] = 14'b0000000_0000000;
		Dminus[5899] = 14'b0000000_0000000;
		Dminus[5900] = 14'b0000000_0000000;
		Dminus[5901] = 14'b0000000_0000000;
		Dminus[5902] = 14'b0000000_0000000;
		Dminus[5903] = 14'b0000000_0000000;
		Dminus[5904] = 14'b0000000_0000000;
		Dminus[5905] = 14'b0000000_0000000;
		Dminus[5906] = 14'b0000000_0000000;
		Dminus[5907] = 14'b0000000_0000000;
		Dminus[5908] = 14'b0000000_0000000;
		Dminus[5909] = 14'b0000000_0000000;
		Dminus[5910] = 14'b0000000_0000000;
		Dminus[5911] = 14'b0000000_0000000;
		Dminus[5912] = 14'b0000000_0000000;
		Dminus[5913] = 14'b0000000_0000000;
		Dminus[5914] = 14'b0000000_0000000;
		Dminus[5915] = 14'b0000000_0000000;
		Dminus[5916] = 14'b0000000_0000000;
		Dminus[5917] = 14'b0000000_0000000;
		Dminus[5918] = 14'b0000000_0000000;
		Dminus[5919] = 14'b0000000_0000000;
		Dminus[5920] = 14'b0000000_0000000;
		Dminus[5921] = 14'b0000000_0000000;
		Dminus[5922] = 14'b0000000_0000000;
		Dminus[5923] = 14'b0000000_0000000;
		Dminus[5924] = 14'b0000000_0000000;
		Dminus[5925] = 14'b0000000_0000000;
		Dminus[5926] = 14'b0000000_0000000;
		Dminus[5927] = 14'b0000000_0000000;
		Dminus[5928] = 14'b0000000_0000000;
		Dminus[5929] = 14'b0000000_0000000;
		Dminus[5930] = 14'b0000000_0000000;
		Dminus[5931] = 14'b0000000_0000000;
		Dminus[5932] = 14'b0000000_0000000;
		Dminus[5933] = 14'b0000000_0000000;
		Dminus[5934] = 14'b0000000_0000000;
		Dminus[5935] = 14'b0000000_0000000;
		Dminus[5936] = 14'b0000000_0000000;
		Dminus[5937] = 14'b0000000_0000000;
		Dminus[5938] = 14'b0000000_0000000;
		Dminus[5939] = 14'b0000000_0000000;
		Dminus[5940] = 14'b0000000_0000000;
		Dminus[5941] = 14'b0000000_0000000;
		Dminus[5942] = 14'b0000000_0000000;
		Dminus[5943] = 14'b0000000_0000000;
		Dminus[5944] = 14'b0000000_0000000;
		Dminus[5945] = 14'b0000000_0000000;
		Dminus[5946] = 14'b0000000_0000000;
		Dminus[5947] = 14'b0000000_0000000;
		Dminus[5948] = 14'b0000000_0000000;
		Dminus[5949] = 14'b0000000_0000000;
		Dminus[5950] = 14'b0000000_0000000;
		Dminus[5951] = 14'b0000000_0000000;
		Dminus[5952] = 14'b0000000_0000000;
		Dminus[5953] = 14'b0000000_0000000;
		Dminus[5954] = 14'b0000000_0000000;
		Dminus[5955] = 14'b0000000_0000000;
		Dminus[5956] = 14'b0000000_0000000;
		Dminus[5957] = 14'b0000000_0000000;
		Dminus[5958] = 14'b0000000_0000000;
		Dminus[5959] = 14'b0000000_0000000;
		Dminus[5960] = 14'b0000000_0000000;
		Dminus[5961] = 14'b0000000_0000000;
		Dminus[5962] = 14'b0000000_0000000;
		Dminus[5963] = 14'b0000000_0000000;
		Dminus[5964] = 14'b0000000_0000000;
		Dminus[5965] = 14'b0000000_0000000;
		Dminus[5966] = 14'b0000000_0000000;
		Dminus[5967] = 14'b0000000_0000000;
		Dminus[5968] = 14'b0000000_0000000;
		Dminus[5969] = 14'b0000000_0000000;
		Dminus[5970] = 14'b0000000_0000000;
		Dminus[5971] = 14'b0000000_0000000;
		Dminus[5972] = 14'b0000000_0000000;
		Dminus[5973] = 14'b0000000_0000000;
		Dminus[5974] = 14'b0000000_0000000;
		Dminus[5975] = 14'b0000000_0000000;
		Dminus[5976] = 14'b0000000_0000000;
		Dminus[5977] = 14'b0000000_0000000;
		Dminus[5978] = 14'b0000000_0000000;
		Dminus[5979] = 14'b0000000_0000000;
		Dminus[5980] = 14'b0000000_0000000;
		Dminus[5981] = 14'b0000000_0000000;
		Dminus[5982] = 14'b0000000_0000000;
		Dminus[5983] = 14'b0000000_0000000;
		Dminus[5984] = 14'b0000000_0000000;
		Dminus[5985] = 14'b0000000_0000000;
		Dminus[5986] = 14'b0000000_0000000;
		Dminus[5987] = 14'b0000000_0000000;
		Dminus[5988] = 14'b0000000_0000000;
		Dminus[5989] = 14'b0000000_0000000;
		Dminus[5990] = 14'b0000000_0000000;
		Dminus[5991] = 14'b0000000_0000000;
		Dminus[5992] = 14'b0000000_0000000;
		Dminus[5993] = 14'b0000000_0000000;
		Dminus[5994] = 14'b0000000_0000000;
		Dminus[5995] = 14'b0000000_0000000;
		Dminus[5996] = 14'b0000000_0000000;
		Dminus[5997] = 14'b0000000_0000000;
		Dminus[5998] = 14'b0000000_0000000;
		Dminus[5999] = 14'b0000000_0000000;
		Dminus[6000] = 14'b0000000_0000000;
		Dminus[6001] = 14'b0000000_0000000;
		Dminus[6002] = 14'b0000000_0000000;
		Dminus[6003] = 14'b0000000_0000000;
		Dminus[6004] = 14'b0000000_0000000;
		Dminus[6005] = 14'b0000000_0000000;
		Dminus[6006] = 14'b0000000_0000000;
		Dminus[6007] = 14'b0000000_0000000;
		Dminus[6008] = 14'b0000000_0000000;
		Dminus[6009] = 14'b0000000_0000000;
		Dminus[6010] = 14'b0000000_0000000;
		Dminus[6011] = 14'b0000000_0000000;
		Dminus[6012] = 14'b0000000_0000000;
		Dminus[6013] = 14'b0000000_0000000;
		Dminus[6014] = 14'b0000000_0000000;
		Dminus[6015] = 14'b0000000_0000000;
		Dminus[6016] = 14'b0000000_0000000;
		Dminus[6017] = 14'b0000000_0000000;
		Dminus[6018] = 14'b0000000_0000000;
		Dminus[6019] = 14'b0000000_0000000;
		Dminus[6020] = 14'b0000000_0000000;
		Dminus[6021] = 14'b0000000_0000000;
		Dminus[6022] = 14'b0000000_0000000;
		Dminus[6023] = 14'b0000000_0000000;
		Dminus[6024] = 14'b0000000_0000000;
		Dminus[6025] = 14'b0000000_0000000;
		Dminus[6026] = 14'b0000000_0000000;
		Dminus[6027] = 14'b0000000_0000000;
		Dminus[6028] = 14'b0000000_0000000;
		Dminus[6029] = 14'b0000000_0000000;
		Dminus[6030] = 14'b0000000_0000000;
		Dminus[6031] = 14'b0000000_0000000;
		Dminus[6032] = 14'b0000000_0000000;
		Dminus[6033] = 14'b0000000_0000000;
		Dminus[6034] = 14'b0000000_0000000;
		Dminus[6035] = 14'b0000000_0000000;
		Dminus[6036] = 14'b0000000_0000000;
		Dminus[6037] = 14'b0000000_0000000;
		Dminus[6038] = 14'b0000000_0000000;
		Dminus[6039] = 14'b0000000_0000000;
		Dminus[6040] = 14'b0000000_0000000;
		Dminus[6041] = 14'b0000000_0000000;
		Dminus[6042] = 14'b0000000_0000000;
		Dminus[6043] = 14'b0000000_0000000;
		Dminus[6044] = 14'b0000000_0000000;
		Dminus[6045] = 14'b0000000_0000000;
		Dminus[6046] = 14'b0000000_0000000;
		Dminus[6047] = 14'b0000000_0000000;
		Dminus[6048] = 14'b0000000_0000000;
		Dminus[6049] = 14'b0000000_0000000;
		Dminus[6050] = 14'b0000000_0000000;
		Dminus[6051] = 14'b0000000_0000000;
		Dminus[6052] = 14'b0000000_0000000;
		Dminus[6053] = 14'b0000000_0000000;
		Dminus[6054] = 14'b0000000_0000000;
		Dminus[6055] = 14'b0000000_0000000;
		Dminus[6056] = 14'b0000000_0000000;
		Dminus[6057] = 14'b0000000_0000000;
		Dminus[6058] = 14'b0000000_0000000;
		Dminus[6059] = 14'b0000000_0000000;
		Dminus[6060] = 14'b0000000_0000000;
		Dminus[6061] = 14'b0000000_0000000;
		Dminus[6062] = 14'b0000000_0000000;
		Dminus[6063] = 14'b0000000_0000000;
		Dminus[6064] = 14'b0000000_0000000;
		Dminus[6065] = 14'b0000000_0000000;
		Dminus[6066] = 14'b0000000_0000000;
		Dminus[6067] = 14'b0000000_0000000;
		Dminus[6068] = 14'b0000000_0000000;
		Dminus[6069] = 14'b0000000_0000000;
		Dminus[6070] = 14'b0000000_0000000;
		Dminus[6071] = 14'b0000000_0000000;
		Dminus[6072] = 14'b0000000_0000000;
		Dminus[6073] = 14'b0000000_0000000;
		Dminus[6074] = 14'b0000000_0000000;
		Dminus[6075] = 14'b0000000_0000000;
		Dminus[6076] = 14'b0000000_0000000;
		Dminus[6077] = 14'b0000000_0000000;
		Dminus[6078] = 14'b0000000_0000000;
		Dminus[6079] = 14'b0000000_0000000;
		Dminus[6080] = 14'b0000000_0000000;
		Dminus[6081] = 14'b0000000_0000000;
		Dminus[6082] = 14'b0000000_0000000;
		Dminus[6083] = 14'b0000000_0000000;
		Dminus[6084] = 14'b0000000_0000000;
		Dminus[6085] = 14'b0000000_0000000;
		Dminus[6086] = 14'b0000000_0000000;
		Dminus[6087] = 14'b0000000_0000000;
		Dminus[6088] = 14'b0000000_0000000;
		Dminus[6089] = 14'b0000000_0000000;
		Dminus[6090] = 14'b0000000_0000000;
		Dminus[6091] = 14'b0000000_0000000;
		Dminus[6092] = 14'b0000000_0000000;
		Dminus[6093] = 14'b0000000_0000000;
		Dminus[6094] = 14'b0000000_0000000;
		Dminus[6095] = 14'b0000000_0000000;
		Dminus[6096] = 14'b0000000_0000000;
		Dminus[6097] = 14'b0000000_0000000;
		Dminus[6098] = 14'b0000000_0000000;
		Dminus[6099] = 14'b0000000_0000000;
		Dminus[6100] = 14'b0000000_0000000;
		Dminus[6101] = 14'b0000000_0000000;
		Dminus[6102] = 14'b0000000_0000000;
		Dminus[6103] = 14'b0000000_0000000;
		Dminus[6104] = 14'b0000000_0000000;
		Dminus[6105] = 14'b0000000_0000000;
		Dminus[6106] = 14'b0000000_0000000;
		Dminus[6107] = 14'b0000000_0000000;
		Dminus[6108] = 14'b0000000_0000000;
		Dminus[6109] = 14'b0000000_0000000;
		Dminus[6110] = 14'b0000000_0000000;
		Dminus[6111] = 14'b0000000_0000000;
		Dminus[6112] = 14'b0000000_0000000;
		Dminus[6113] = 14'b0000000_0000000;
		Dminus[6114] = 14'b0000000_0000000;
		Dminus[6115] = 14'b0000000_0000000;
		Dminus[6116] = 14'b0000000_0000000;
		Dminus[6117] = 14'b0000000_0000000;
		Dminus[6118] = 14'b0000000_0000000;
		Dminus[6119] = 14'b0000000_0000000;
		Dminus[6120] = 14'b0000000_0000000;
		Dminus[6121] = 14'b0000000_0000000;
		Dminus[6122] = 14'b0000000_0000000;
		Dminus[6123] = 14'b0000000_0000000;
		Dminus[6124] = 14'b0000000_0000000;
		Dminus[6125] = 14'b0000000_0000000;
		Dminus[6126] = 14'b0000000_0000000;
		Dminus[6127] = 14'b0000000_0000000;
		Dminus[6128] = 14'b0000000_0000000;
		Dminus[6129] = 14'b0000000_0000000;
		Dminus[6130] = 14'b0000000_0000000;
		Dminus[6131] = 14'b0000000_0000000;
		Dminus[6132] = 14'b0000000_0000000;
		Dminus[6133] = 14'b0000000_0000000;
		Dminus[6134] = 14'b0000000_0000000;
		Dminus[6135] = 14'b0000000_0000000;
		Dminus[6136] = 14'b0000000_0000000;
		Dminus[6137] = 14'b0000000_0000000;
		Dminus[6138] = 14'b0000000_0000000;
		Dminus[6139] = 14'b0000000_0000000;
		Dminus[6140] = 14'b0000000_0000000;
		Dminus[6141] = 14'b0000000_0000000;
		Dminus[6142] = 14'b0000000_0000000;
		Dminus[6143] = 14'b0000000_0000000;
		Dminus[6144] = 14'b0000000_0000000;
		Dminus[6145] = 14'b0000000_0000000;
		Dminus[6146] = 14'b0000000_0000000;
		Dminus[6147] = 14'b0000000_0000000;
		Dminus[6148] = 14'b0000000_0000000;
		Dminus[6149] = 14'b0000000_0000000;
		Dminus[6150] = 14'b0000000_0000000;
		Dminus[6151] = 14'b0000000_0000000;
		Dminus[6152] = 14'b0000000_0000000;
		Dminus[6153] = 14'b0000000_0000000;
		Dminus[6154] = 14'b0000000_0000000;
		Dminus[6155] = 14'b0000000_0000000;
		Dminus[6156] = 14'b0000000_0000000;
		Dminus[6157] = 14'b0000000_0000000;
		Dminus[6158] = 14'b0000000_0000000;
		Dminus[6159] = 14'b0000000_0000000;
		Dminus[6160] = 14'b0000000_0000000;
		Dminus[6161] = 14'b0000000_0000000;
		Dminus[6162] = 14'b0000000_0000000;
		Dminus[6163] = 14'b0000000_0000000;
		Dminus[6164] = 14'b0000000_0000000;
		Dminus[6165] = 14'b0000000_0000000;
		Dminus[6166] = 14'b0000000_0000000;
		Dminus[6167] = 14'b0000000_0000000;
		Dminus[6168] = 14'b0000000_0000000;
		Dminus[6169] = 14'b0000000_0000000;
		Dminus[6170] = 14'b0000000_0000000;
		Dminus[6171] = 14'b0000000_0000000;
		Dminus[6172] = 14'b0000000_0000000;
		Dminus[6173] = 14'b0000000_0000000;
		Dminus[6174] = 14'b0000000_0000000;
		Dminus[6175] = 14'b0000000_0000000;
		Dminus[6176] = 14'b0000000_0000000;
		Dminus[6177] = 14'b0000000_0000000;
		Dminus[6178] = 14'b0000000_0000000;
		Dminus[6179] = 14'b0000000_0000000;
		Dminus[6180] = 14'b0000000_0000000;
		Dminus[6181] = 14'b0000000_0000000;
		Dminus[6182] = 14'b0000000_0000000;
		Dminus[6183] = 14'b0000000_0000000;
		Dminus[6184] = 14'b0000000_0000000;
		Dminus[6185] = 14'b0000000_0000000;
		Dminus[6186] = 14'b0000000_0000000;
		Dminus[6187] = 14'b0000000_0000000;
		Dminus[6188] = 14'b0000000_0000000;
		Dminus[6189] = 14'b0000000_0000000;
		Dminus[6190] = 14'b0000000_0000000;
		Dminus[6191] = 14'b0000000_0000000;
		Dminus[6192] = 14'b0000000_0000000;
		Dminus[6193] = 14'b0000000_0000000;
		Dminus[6194] = 14'b0000000_0000000;
		Dminus[6195] = 14'b0000000_0000000;
		Dminus[6196] = 14'b0000000_0000000;
		Dminus[6197] = 14'b0000000_0000000;
		Dminus[6198] = 14'b0000000_0000000;
		Dminus[6199] = 14'b0000000_0000000;
		Dminus[6200] = 14'b0000000_0000000;
		Dminus[6201] = 14'b0000000_0000000;
		Dminus[6202] = 14'b0000000_0000000;
		Dminus[6203] = 14'b0000000_0000000;
		Dminus[6204] = 14'b0000000_0000000;
		Dminus[6205] = 14'b0000000_0000000;
		Dminus[6206] = 14'b0000000_0000000;
		Dminus[6207] = 14'b0000000_0000000;
		Dminus[6208] = 14'b0000000_0000000;
		Dminus[6209] = 14'b0000000_0000000;
		Dminus[6210] = 14'b0000000_0000000;
		Dminus[6211] = 14'b0000000_0000000;
		Dminus[6212] = 14'b0000000_0000000;
		Dminus[6213] = 14'b0000000_0000000;
		Dminus[6214] = 14'b0000000_0000000;
		Dminus[6215] = 14'b0000000_0000000;
		Dminus[6216] = 14'b0000000_0000000;
		Dminus[6217] = 14'b0000000_0000000;
		Dminus[6218] = 14'b0000000_0000000;
		Dminus[6219] = 14'b0000000_0000000;
		Dminus[6220] = 14'b0000000_0000000;
		Dminus[6221] = 14'b0000000_0000000;
		Dminus[6222] = 14'b0000000_0000000;
		Dminus[6223] = 14'b0000000_0000000;
		Dminus[6224] = 14'b0000000_0000000;
		Dminus[6225] = 14'b0000000_0000000;
		Dminus[6226] = 14'b0000000_0000000;
		Dminus[6227] = 14'b0000000_0000000;
		Dminus[6228] = 14'b0000000_0000000;
		Dminus[6229] = 14'b0000000_0000000;
		Dminus[6230] = 14'b0000000_0000000;
		Dminus[6231] = 14'b0000000_0000000;
		Dminus[6232] = 14'b0000000_0000000;
		Dminus[6233] = 14'b0000000_0000000;
		Dminus[6234] = 14'b0000000_0000000;
		Dminus[6235] = 14'b0000000_0000000;
		Dminus[6236] = 14'b0000000_0000000;
		Dminus[6237] = 14'b0000000_0000000;
		Dminus[6238] = 14'b0000000_0000000;
		Dminus[6239] = 14'b0000000_0000000;
		Dminus[6240] = 14'b0000000_0000000;
		Dminus[6241] = 14'b0000000_0000000;
		Dminus[6242] = 14'b0000000_0000000;
		Dminus[6243] = 14'b0000000_0000000;
		Dminus[6244] = 14'b0000000_0000000;
		Dminus[6245] = 14'b0000000_0000000;
		Dminus[6246] = 14'b0000000_0000000;
		Dminus[6247] = 14'b0000000_0000000;
		Dminus[6248] = 14'b0000000_0000000;
		Dminus[6249] = 14'b0000000_0000000;
		Dminus[6250] = 14'b0000000_0000000;
		Dminus[6251] = 14'b0000000_0000000;
		Dminus[6252] = 14'b0000000_0000000;
		Dminus[6253] = 14'b0000000_0000000;
		Dminus[6254] = 14'b0000000_0000000;
		Dminus[6255] = 14'b0000000_0000000;
		Dminus[6256] = 14'b0000000_0000000;
		Dminus[6257] = 14'b0000000_0000000;
		Dminus[6258] = 14'b0000000_0000000;
		Dminus[6259] = 14'b0000000_0000000;
		Dminus[6260] = 14'b0000000_0000000;
		Dminus[6261] = 14'b0000000_0000000;
		Dminus[6262] = 14'b0000000_0000000;
		Dminus[6263] = 14'b0000000_0000000;
		Dminus[6264] = 14'b0000000_0000000;
		Dminus[6265] = 14'b0000000_0000000;
		Dminus[6266] = 14'b0000000_0000000;
		Dminus[6267] = 14'b0000000_0000000;
		Dminus[6268] = 14'b0000000_0000000;
		Dminus[6269] = 14'b0000000_0000000;
		Dminus[6270] = 14'b0000000_0000000;
		Dminus[6271] = 14'b0000000_0000000;
		Dminus[6272] = 14'b0000000_0000000;
		Dminus[6273] = 14'b0000000_0000000;
		Dminus[6274] = 14'b0000000_0000000;
		Dminus[6275] = 14'b0000000_0000000;
		Dminus[6276] = 14'b0000000_0000000;
		Dminus[6277] = 14'b0000000_0000000;
		Dminus[6278] = 14'b0000000_0000000;
		Dminus[6279] = 14'b0000000_0000000;
		Dminus[6280] = 14'b0000000_0000000;
		Dminus[6281] = 14'b0000000_0000000;
		Dminus[6282] = 14'b0000000_0000000;
		Dminus[6283] = 14'b0000000_0000000;
		Dminus[6284] = 14'b0000000_0000000;
		Dminus[6285] = 14'b0000000_0000000;
		Dminus[6286] = 14'b0000000_0000000;
		Dminus[6287] = 14'b0000000_0000000;
		Dminus[6288] = 14'b0000000_0000000;
		Dminus[6289] = 14'b0000000_0000000;
		Dminus[6290] = 14'b0000000_0000000;
		Dminus[6291] = 14'b0000000_0000000;
		Dminus[6292] = 14'b0000000_0000000;
		Dminus[6293] = 14'b0000000_0000000;
		Dminus[6294] = 14'b0000000_0000000;
		Dminus[6295] = 14'b0000000_0000000;
		Dminus[6296] = 14'b0000000_0000000;
		Dminus[6297] = 14'b0000000_0000000;
		Dminus[6298] = 14'b0000000_0000000;
		Dminus[6299] = 14'b0000000_0000000;
		Dminus[6300] = 14'b0000000_0000000;
		Dminus[6301] = 14'b0000000_0000000;
		Dminus[6302] = 14'b0000000_0000000;
		Dminus[6303] = 14'b0000000_0000000;
		Dminus[6304] = 14'b0000000_0000000;
		Dminus[6305] = 14'b0000000_0000000;
		Dminus[6306] = 14'b0000000_0000000;
		Dminus[6307] = 14'b0000000_0000000;
		Dminus[6308] = 14'b0000000_0000000;
		Dminus[6309] = 14'b0000000_0000000;
		Dminus[6310] = 14'b0000000_0000000;
		Dminus[6311] = 14'b0000000_0000000;
		Dminus[6312] = 14'b0000000_0000000;
		Dminus[6313] = 14'b0000000_0000000;
		Dminus[6314] = 14'b0000000_0000000;
		Dminus[6315] = 14'b0000000_0000000;
		Dminus[6316] = 14'b0000000_0000000;
		Dminus[6317] = 14'b0000000_0000000;
		Dminus[6318] = 14'b0000000_0000000;
		Dminus[6319] = 14'b0000000_0000000;
		Dminus[6320] = 14'b0000000_0000000;
		Dminus[6321] = 14'b0000000_0000000;
		Dminus[6322] = 14'b0000000_0000000;
		Dminus[6323] = 14'b0000000_0000000;
		Dminus[6324] = 14'b0000000_0000000;
		Dminus[6325] = 14'b0000000_0000000;
		Dminus[6326] = 14'b0000000_0000000;
		Dminus[6327] = 14'b0000000_0000000;
		Dminus[6328] = 14'b0000000_0000000;
		Dminus[6329] = 14'b0000000_0000000;
		Dminus[6330] = 14'b0000000_0000000;
		Dminus[6331] = 14'b0000000_0000000;
		Dminus[6332] = 14'b0000000_0000000;
		Dminus[6333] = 14'b0000000_0000000;
		Dminus[6334] = 14'b0000000_0000000;
		Dminus[6335] = 14'b0000000_0000000;
		Dminus[6336] = 14'b0000000_0000000;
		Dminus[6337] = 14'b0000000_0000000;
		Dminus[6338] = 14'b0000000_0000000;
		Dminus[6339] = 14'b0000000_0000000;
		Dminus[6340] = 14'b0000000_0000000;
		Dminus[6341] = 14'b0000000_0000000;
		Dminus[6342] = 14'b0000000_0000000;
		Dminus[6343] = 14'b0000000_0000000;
		Dminus[6344] = 14'b0000000_0000000;
		Dminus[6345] = 14'b0000000_0000000;
		Dminus[6346] = 14'b0000000_0000000;
		Dminus[6347] = 14'b0000000_0000000;
		Dminus[6348] = 14'b0000000_0000000;
		Dminus[6349] = 14'b0000000_0000000;
		Dminus[6350] = 14'b0000000_0000000;
		Dminus[6351] = 14'b0000000_0000000;
		Dminus[6352] = 14'b0000000_0000000;
		Dminus[6353] = 14'b0000000_0000000;
		Dminus[6354] = 14'b0000000_0000000;
		Dminus[6355] = 14'b0000000_0000000;
		Dminus[6356] = 14'b0000000_0000000;
		Dminus[6357] = 14'b0000000_0000000;
		Dminus[6358] = 14'b0000000_0000000;
		Dminus[6359] = 14'b0000000_0000000;
		Dminus[6360] = 14'b0000000_0000000;
		Dminus[6361] = 14'b0000000_0000000;
		Dminus[6362] = 14'b0000000_0000000;
		Dminus[6363] = 14'b0000000_0000000;
		Dminus[6364] = 14'b0000000_0000000;
		Dminus[6365] = 14'b0000000_0000000;
		Dminus[6366] = 14'b0000000_0000000;
		Dminus[6367] = 14'b0000000_0000000;
		Dminus[6368] = 14'b0000000_0000000;
		Dminus[6369] = 14'b0000000_0000000;
		Dminus[6370] = 14'b0000000_0000000;
		Dminus[6371] = 14'b0000000_0000000;
		Dminus[6372] = 14'b0000000_0000000;
		Dminus[6373] = 14'b0000000_0000000;
		Dminus[6374] = 14'b0000000_0000000;
		Dminus[6375] = 14'b0000000_0000000;
		Dminus[6376] = 14'b0000000_0000000;
		Dminus[6377] = 14'b0000000_0000000;
		Dminus[6378] = 14'b0000000_0000000;
		Dminus[6379] = 14'b0000000_0000000;
		Dminus[6380] = 14'b0000000_0000000;
		Dminus[6381] = 14'b0000000_0000000;
		Dminus[6382] = 14'b0000000_0000000;
		Dminus[6383] = 14'b0000000_0000000;
		Dminus[6384] = 14'b0000000_0000000;
		Dminus[6385] = 14'b0000000_0000000;
		Dminus[6386] = 14'b0000000_0000000;
		Dminus[6387] = 14'b0000000_0000000;
		Dminus[6388] = 14'b0000000_0000000;
		Dminus[6389] = 14'b0000000_0000000;
		Dminus[6390] = 14'b0000000_0000000;
		Dminus[6391] = 14'b0000000_0000000;
		Dminus[6392] = 14'b0000000_0000000;
		Dminus[6393] = 14'b0000000_0000000;
		Dminus[6394] = 14'b0000000_0000000;
		Dminus[6395] = 14'b0000000_0000000;
		Dminus[6396] = 14'b0000000_0000000;
		Dminus[6397] = 14'b0000000_0000000;
		Dminus[6398] = 14'b0000000_0000000;
		Dminus[6399] = 14'b0000000_0000000;
		Dminus[6400] = 14'b0000000_0000000;
		Dminus[6401] = 14'b0000000_0000000;
		Dminus[6402] = 14'b0000000_0000000;
		Dminus[6403] = 14'b0000000_0000000;
		Dminus[6404] = 14'b0000000_0000000;
		Dminus[6405] = 14'b0000000_0000000;
		Dminus[6406] = 14'b0000000_0000000;
		Dminus[6407] = 14'b0000000_0000000;
		Dminus[6408] = 14'b0000000_0000000;
		Dminus[6409] = 14'b0000000_0000000;
		Dminus[6410] = 14'b0000000_0000000;
		Dminus[6411] = 14'b0000000_0000000;
		Dminus[6412] = 14'b0000000_0000000;
		Dminus[6413] = 14'b0000000_0000000;
		Dminus[6414] = 14'b0000000_0000000;
		Dminus[6415] = 14'b0000000_0000000;
		Dminus[6416] = 14'b0000000_0000000;
		Dminus[6417] = 14'b0000000_0000000;
		Dminus[6418] = 14'b0000000_0000000;
		Dminus[6419] = 14'b0000000_0000000;
		Dminus[6420] = 14'b0000000_0000000;
		Dminus[6421] = 14'b0000000_0000000;
		Dminus[6422] = 14'b0000000_0000000;
		Dminus[6423] = 14'b0000000_0000000;
		Dminus[6424] = 14'b0000000_0000000;
		Dminus[6425] = 14'b0000000_0000000;
		Dminus[6426] = 14'b0000000_0000000;
		Dminus[6427] = 14'b0000000_0000000;
		Dminus[6428] = 14'b0000000_0000000;
		Dminus[6429] = 14'b0000000_0000000;
		Dminus[6430] = 14'b0000000_0000000;
		Dminus[6431] = 14'b0000000_0000000;
		Dminus[6432] = 14'b0000000_0000000;
		Dminus[6433] = 14'b0000000_0000000;
		Dminus[6434] = 14'b0000000_0000000;
		Dminus[6435] = 14'b0000000_0000000;
		Dminus[6436] = 14'b0000000_0000000;
		Dminus[6437] = 14'b0000000_0000000;
		Dminus[6438] = 14'b0000000_0000000;
		Dminus[6439] = 14'b0000000_0000000;
		Dminus[6440] = 14'b0000000_0000000;
		Dminus[6441] = 14'b0000000_0000000;
		Dminus[6442] = 14'b0000000_0000000;
		Dminus[6443] = 14'b0000000_0000000;
		Dminus[6444] = 14'b0000000_0000000;
		Dminus[6445] = 14'b0000000_0000000;
		Dminus[6446] = 14'b0000000_0000000;
		Dminus[6447] = 14'b0000000_0000000;
		Dminus[6448] = 14'b0000000_0000000;
		Dminus[6449] = 14'b0000000_0000000;
		Dminus[6450] = 14'b0000000_0000000;
		Dminus[6451] = 14'b0000000_0000000;
		Dminus[6452] = 14'b0000000_0000000;
		Dminus[6453] = 14'b0000000_0000000;
		Dminus[6454] = 14'b0000000_0000000;
		Dminus[6455] = 14'b0000000_0000000;
		Dminus[6456] = 14'b0000000_0000000;
		Dminus[6457] = 14'b0000000_0000000;
		Dminus[6458] = 14'b0000000_0000000;
		Dminus[6459] = 14'b0000000_0000000;
		Dminus[6460] = 14'b0000000_0000000;
		Dminus[6461] = 14'b0000000_0000000;
		Dminus[6462] = 14'b0000000_0000000;
		Dminus[6463] = 14'b0000000_0000000;
		Dminus[6464] = 14'b0000000_0000000;
		Dminus[6465] = 14'b0000000_0000000;
		Dminus[6466] = 14'b0000000_0000000;
		Dminus[6467] = 14'b0000000_0000000;
		Dminus[6468] = 14'b0000000_0000000;
		Dminus[6469] = 14'b0000000_0000000;
		Dminus[6470] = 14'b0000000_0000000;
		Dminus[6471] = 14'b0000000_0000000;
		Dminus[6472] = 14'b0000000_0000000;
		Dminus[6473] = 14'b0000000_0000000;
		Dminus[6474] = 14'b0000000_0000000;
		Dminus[6475] = 14'b0000000_0000000;
		Dminus[6476] = 14'b0000000_0000000;
		Dminus[6477] = 14'b0000000_0000000;
		Dminus[6478] = 14'b0000000_0000000;
		Dminus[6479] = 14'b0000000_0000000;
		Dminus[6480] = 14'b0000000_0000000;
		Dminus[6481] = 14'b0000000_0000000;
		Dminus[6482] = 14'b0000000_0000000;
		Dminus[6483] = 14'b0000000_0000000;
		Dminus[6484] = 14'b0000000_0000000;
		Dminus[6485] = 14'b0000000_0000000;
		Dminus[6486] = 14'b0000000_0000000;
		Dminus[6487] = 14'b0000000_0000000;
		Dminus[6488] = 14'b0000000_0000000;
		Dminus[6489] = 14'b0000000_0000000;
		Dminus[6490] = 14'b0000000_0000000;
		Dminus[6491] = 14'b0000000_0000000;
		Dminus[6492] = 14'b0000000_0000000;
		Dminus[6493] = 14'b0000000_0000000;
		Dminus[6494] = 14'b0000000_0000000;
		Dminus[6495] = 14'b0000000_0000000;
		Dminus[6496] = 14'b0000000_0000000;
		Dminus[6497] = 14'b0000000_0000000;
		Dminus[6498] = 14'b0000000_0000000;
		Dminus[6499] = 14'b0000000_0000000;
		Dminus[6500] = 14'b0000000_0000000;
		Dminus[6501] = 14'b0000000_0000000;
		Dminus[6502] = 14'b0000000_0000000;
		Dminus[6503] = 14'b0000000_0000000;
		Dminus[6504] = 14'b0000000_0000000;
		Dminus[6505] = 14'b0000000_0000000;
		Dminus[6506] = 14'b0000000_0000000;
		Dminus[6507] = 14'b0000000_0000000;
		Dminus[6508] = 14'b0000000_0000000;
		Dminus[6509] = 14'b0000000_0000000;
		Dminus[6510] = 14'b0000000_0000000;
		Dminus[6511] = 14'b0000000_0000000;
		Dminus[6512] = 14'b0000000_0000000;
		Dminus[6513] = 14'b0000000_0000000;
		Dminus[6514] = 14'b0000000_0000000;
		Dminus[6515] = 14'b0000000_0000000;
		Dminus[6516] = 14'b0000000_0000000;
		Dminus[6517] = 14'b0000000_0000000;
		Dminus[6518] = 14'b0000000_0000000;
		Dminus[6519] = 14'b0000000_0000000;
		Dminus[6520] = 14'b0000000_0000000;
		Dminus[6521] = 14'b0000000_0000000;
		Dminus[6522] = 14'b0000000_0000000;
		Dminus[6523] = 14'b0000000_0000000;
		Dminus[6524] = 14'b0000000_0000000;
		Dminus[6525] = 14'b0000000_0000000;
		Dminus[6526] = 14'b0000000_0000000;
		Dminus[6527] = 14'b0000000_0000000;
		Dminus[6528] = 14'b0000000_0000000;
		Dminus[6529] = 14'b0000000_0000000;
		Dminus[6530] = 14'b0000000_0000000;
		Dminus[6531] = 14'b0000000_0000000;
		Dminus[6532] = 14'b0000000_0000000;
		Dminus[6533] = 14'b0000000_0000000;
		Dminus[6534] = 14'b0000000_0000000;
		Dminus[6535] = 14'b0000000_0000000;
		Dminus[6536] = 14'b0000000_0000000;
		Dminus[6537] = 14'b0000000_0000000;
		Dminus[6538] = 14'b0000000_0000000;
		Dminus[6539] = 14'b0000000_0000000;
		Dminus[6540] = 14'b0000000_0000000;
		Dminus[6541] = 14'b0000000_0000000;
		Dminus[6542] = 14'b0000000_0000000;
		Dminus[6543] = 14'b0000000_0000000;
		Dminus[6544] = 14'b0000000_0000000;
		Dminus[6545] = 14'b0000000_0000000;
		Dminus[6546] = 14'b0000000_0000000;
		Dminus[6547] = 14'b0000000_0000000;
		Dminus[6548] = 14'b0000000_0000000;
		Dminus[6549] = 14'b0000000_0000000;
		Dminus[6550] = 14'b0000000_0000000;
		Dminus[6551] = 14'b0000000_0000000;
		Dminus[6552] = 14'b0000000_0000000;
		Dminus[6553] = 14'b0000000_0000000;
		Dminus[6554] = 14'b0000000_0000000;
		Dminus[6555] = 14'b0000000_0000000;
		Dminus[6556] = 14'b0000000_0000000;
		Dminus[6557] = 14'b0000000_0000000;
		Dminus[6558] = 14'b0000000_0000000;
		Dminus[6559] = 14'b0000000_0000000;
		Dminus[6560] = 14'b0000000_0000000;
		Dminus[6561] = 14'b0000000_0000000;
		Dminus[6562] = 14'b0000000_0000000;
		Dminus[6563] = 14'b0000000_0000000;
		Dminus[6564] = 14'b0000000_0000000;
		Dminus[6565] = 14'b0000000_0000000;
		Dminus[6566] = 14'b0000000_0000000;
		Dminus[6567] = 14'b0000000_0000000;
		Dminus[6568] = 14'b0000000_0000000;
		Dminus[6569] = 14'b0000000_0000000;
		Dminus[6570] = 14'b0000000_0000000;
		Dminus[6571] = 14'b0000000_0000000;
		Dminus[6572] = 14'b0000000_0000000;
		Dminus[6573] = 14'b0000000_0000000;
		Dminus[6574] = 14'b0000000_0000000;
		Dminus[6575] = 14'b0000000_0000000;
		Dminus[6576] = 14'b0000000_0000000;
		Dminus[6577] = 14'b0000000_0000000;
		Dminus[6578] = 14'b0000000_0000000;
		Dminus[6579] = 14'b0000000_0000000;
		Dminus[6580] = 14'b0000000_0000000;
		Dminus[6581] = 14'b0000000_0000000;
		Dminus[6582] = 14'b0000000_0000000;
		Dminus[6583] = 14'b0000000_0000000;
		Dminus[6584] = 14'b0000000_0000000;
		Dminus[6585] = 14'b0000000_0000000;
		Dminus[6586] = 14'b0000000_0000000;
		Dminus[6587] = 14'b0000000_0000000;
		Dminus[6588] = 14'b0000000_0000000;
		Dminus[6589] = 14'b0000000_0000000;
		Dminus[6590] = 14'b0000000_0000000;
		Dminus[6591] = 14'b0000000_0000000;
		Dminus[6592] = 14'b0000000_0000000;
		Dminus[6593] = 14'b0000000_0000000;
		Dminus[6594] = 14'b0000000_0000000;
		Dminus[6595] = 14'b0000000_0000000;
		Dminus[6596] = 14'b0000000_0000000;
		Dminus[6597] = 14'b0000000_0000000;
		Dminus[6598] = 14'b0000000_0000000;
		Dminus[6599] = 14'b0000000_0000000;
		Dminus[6600] = 14'b0000000_0000000;
		Dminus[6601] = 14'b0000000_0000000;
		Dminus[6602] = 14'b0000000_0000000;
		Dminus[6603] = 14'b0000000_0000000;
		Dminus[6604] = 14'b0000000_0000000;
		Dminus[6605] = 14'b0000000_0000000;
		Dminus[6606] = 14'b0000000_0000000;
		Dminus[6607] = 14'b0000000_0000000;
		Dminus[6608] = 14'b0000000_0000000;
		Dminus[6609] = 14'b0000000_0000000;
		Dminus[6610] = 14'b0000000_0000000;
		Dminus[6611] = 14'b0000000_0000000;
		Dminus[6612] = 14'b0000000_0000000;
		Dminus[6613] = 14'b0000000_0000000;
		Dminus[6614] = 14'b0000000_0000000;
		Dminus[6615] = 14'b0000000_0000000;
		Dminus[6616] = 14'b0000000_0000000;
		Dminus[6617] = 14'b0000000_0000000;
		Dminus[6618] = 14'b0000000_0000000;
		Dminus[6619] = 14'b0000000_0000000;
		Dminus[6620] = 14'b0000000_0000000;
		Dminus[6621] = 14'b0000000_0000000;
		Dminus[6622] = 14'b0000000_0000000;
		Dminus[6623] = 14'b0000000_0000000;
		Dminus[6624] = 14'b0000000_0000000;
		Dminus[6625] = 14'b0000000_0000000;
		Dminus[6626] = 14'b0000000_0000000;
		Dminus[6627] = 14'b0000000_0000000;
		Dminus[6628] = 14'b0000000_0000000;
		Dminus[6629] = 14'b0000000_0000000;
		Dminus[6630] = 14'b0000000_0000000;
		Dminus[6631] = 14'b0000000_0000000;
		Dminus[6632] = 14'b0000000_0000000;
		Dminus[6633] = 14'b0000000_0000000;
		Dminus[6634] = 14'b0000000_0000000;
		Dminus[6635] = 14'b0000000_0000000;
		Dminus[6636] = 14'b0000000_0000000;
		Dminus[6637] = 14'b0000000_0000000;
		Dminus[6638] = 14'b0000000_0000000;
		Dminus[6639] = 14'b0000000_0000000;
		Dminus[6640] = 14'b0000000_0000000;
		Dminus[6641] = 14'b0000000_0000000;
		Dminus[6642] = 14'b0000000_0000000;
		Dminus[6643] = 14'b0000000_0000000;
		Dminus[6644] = 14'b0000000_0000000;
		Dminus[6645] = 14'b0000000_0000000;
		Dminus[6646] = 14'b0000000_0000000;
		Dminus[6647] = 14'b0000000_0000000;
		Dminus[6648] = 14'b0000000_0000000;
		Dminus[6649] = 14'b0000000_0000000;
		Dminus[6650] = 14'b0000000_0000000;
		Dminus[6651] = 14'b0000000_0000000;
		Dminus[6652] = 14'b0000000_0000000;
		Dminus[6653] = 14'b0000000_0000000;
		Dminus[6654] = 14'b0000000_0000000;
		Dminus[6655] = 14'b0000000_0000000;
		Dminus[6656] = 14'b0000000_0000000;
		Dminus[6657] = 14'b0000000_0000000;
		Dminus[6658] = 14'b0000000_0000000;
		Dminus[6659] = 14'b0000000_0000000;
		Dminus[6660] = 14'b0000000_0000000;
		Dminus[6661] = 14'b0000000_0000000;
		Dminus[6662] = 14'b0000000_0000000;
		Dminus[6663] = 14'b0000000_0000000;
		Dminus[6664] = 14'b0000000_0000000;
		Dminus[6665] = 14'b0000000_0000000;
		Dminus[6666] = 14'b0000000_0000000;
		Dminus[6667] = 14'b0000000_0000000;
		Dminus[6668] = 14'b0000000_0000000;
		Dminus[6669] = 14'b0000000_0000000;
		Dminus[6670] = 14'b0000000_0000000;
		Dminus[6671] = 14'b0000000_0000000;
		Dminus[6672] = 14'b0000000_0000000;
		Dminus[6673] = 14'b0000000_0000000;
		Dminus[6674] = 14'b0000000_0000000;
		Dminus[6675] = 14'b0000000_0000000;
		Dminus[6676] = 14'b0000000_0000000;
		Dminus[6677] = 14'b0000000_0000000;
		Dminus[6678] = 14'b0000000_0000000;
		Dminus[6679] = 14'b0000000_0000000;
		Dminus[6680] = 14'b0000000_0000000;
		Dminus[6681] = 14'b0000000_0000000;
		Dminus[6682] = 14'b0000000_0000000;
		Dminus[6683] = 14'b0000000_0000000;
		Dminus[6684] = 14'b0000000_0000000;
		Dminus[6685] = 14'b0000000_0000000;
		Dminus[6686] = 14'b0000000_0000000;
		Dminus[6687] = 14'b0000000_0000000;
		Dminus[6688] = 14'b0000000_0000000;
		Dminus[6689] = 14'b0000000_0000000;
		Dminus[6690] = 14'b0000000_0000000;
		Dminus[6691] = 14'b0000000_0000000;
		Dminus[6692] = 14'b0000000_0000000;
		Dminus[6693] = 14'b0000000_0000000;
		Dminus[6694] = 14'b0000000_0000000;
		Dminus[6695] = 14'b0000000_0000000;
		Dminus[6696] = 14'b0000000_0000000;
		Dminus[6697] = 14'b0000000_0000000;
		Dminus[6698] = 14'b0000000_0000000;
		Dminus[6699] = 14'b0000000_0000000;
		Dminus[6700] = 14'b0000000_0000000;
		Dminus[6701] = 14'b0000000_0000000;
		Dminus[6702] = 14'b0000000_0000000;
		Dminus[6703] = 14'b0000000_0000000;
		Dminus[6704] = 14'b0000000_0000000;
		Dminus[6705] = 14'b0000000_0000000;
		Dminus[6706] = 14'b0000000_0000000;
		Dminus[6707] = 14'b0000000_0000000;
		Dminus[6708] = 14'b0000000_0000000;
		Dminus[6709] = 14'b0000000_0000000;
		Dminus[6710] = 14'b0000000_0000000;
		Dminus[6711] = 14'b0000000_0000000;
		Dminus[6712] = 14'b0000000_0000000;
		Dminus[6713] = 14'b0000000_0000000;
		Dminus[6714] = 14'b0000000_0000000;
		Dminus[6715] = 14'b0000000_0000000;
		Dminus[6716] = 14'b0000000_0000000;
		Dminus[6717] = 14'b0000000_0000000;
		Dminus[6718] = 14'b0000000_0000000;
		Dminus[6719] = 14'b0000000_0000000;
		Dminus[6720] = 14'b0000000_0000000;
		Dminus[6721] = 14'b0000000_0000000;
		Dminus[6722] = 14'b0000000_0000000;
		Dminus[6723] = 14'b0000000_0000000;
		Dminus[6724] = 14'b0000000_0000000;
		Dminus[6725] = 14'b0000000_0000000;
		Dminus[6726] = 14'b0000000_0000000;
		Dminus[6727] = 14'b0000000_0000000;
		Dminus[6728] = 14'b0000000_0000000;
		Dminus[6729] = 14'b0000000_0000000;
		Dminus[6730] = 14'b0000000_0000000;
		Dminus[6731] = 14'b0000000_0000000;
		Dminus[6732] = 14'b0000000_0000000;
		Dminus[6733] = 14'b0000000_0000000;
		Dminus[6734] = 14'b0000000_0000000;
		Dminus[6735] = 14'b0000000_0000000;
		Dminus[6736] = 14'b0000000_0000000;
		Dminus[6737] = 14'b0000000_0000000;
		Dminus[6738] = 14'b0000000_0000000;
		Dminus[6739] = 14'b0000000_0000000;
		Dminus[6740] = 14'b0000000_0000000;
		Dminus[6741] = 14'b0000000_0000000;
		Dminus[6742] = 14'b0000000_0000000;
		Dminus[6743] = 14'b0000000_0000000;
		Dminus[6744] = 14'b0000000_0000000;
		Dminus[6745] = 14'b0000000_0000000;
		Dminus[6746] = 14'b0000000_0000000;
		Dminus[6747] = 14'b0000000_0000000;
		Dminus[6748] = 14'b0000000_0000000;
		Dminus[6749] = 14'b0000000_0000000;
		Dminus[6750] = 14'b0000000_0000000;
		Dminus[6751] = 14'b0000000_0000000;
		Dminus[6752] = 14'b0000000_0000000;
		Dminus[6753] = 14'b0000000_0000000;
		Dminus[6754] = 14'b0000000_0000000;
		Dminus[6755] = 14'b0000000_0000000;
		Dminus[6756] = 14'b0000000_0000000;
		Dminus[6757] = 14'b0000000_0000000;
		Dminus[6758] = 14'b0000000_0000000;
		Dminus[6759] = 14'b0000000_0000000;
		Dminus[6760] = 14'b0000000_0000000;
		Dminus[6761] = 14'b0000000_0000000;
		Dminus[6762] = 14'b0000000_0000000;
		Dminus[6763] = 14'b0000000_0000000;
		Dminus[6764] = 14'b0000000_0000000;
		Dminus[6765] = 14'b0000000_0000000;
		Dminus[6766] = 14'b0000000_0000000;
		Dminus[6767] = 14'b0000000_0000000;
		Dminus[6768] = 14'b0000000_0000000;
		Dminus[6769] = 14'b0000000_0000000;
		Dminus[6770] = 14'b0000000_0000000;
		Dminus[6771] = 14'b0000000_0000000;
		Dminus[6772] = 14'b0000000_0000000;
		Dminus[6773] = 14'b0000000_0000000;
		Dminus[6774] = 14'b0000000_0000000;
		Dminus[6775] = 14'b0000000_0000000;
		Dminus[6776] = 14'b0000000_0000000;
		Dminus[6777] = 14'b0000000_0000000;
		Dminus[6778] = 14'b0000000_0000000;
		Dminus[6779] = 14'b0000000_0000000;
		Dminus[6780] = 14'b0000000_0000000;
		Dminus[6781] = 14'b0000000_0000000;
		Dminus[6782] = 14'b0000000_0000000;
		Dminus[6783] = 14'b0000000_0000000;
		Dminus[6784] = 14'b0000000_0000000;
		Dminus[6785] = 14'b0000000_0000000;
		Dminus[6786] = 14'b0000000_0000000;
		Dminus[6787] = 14'b0000000_0000000;
		Dminus[6788] = 14'b0000000_0000000;
		Dminus[6789] = 14'b0000000_0000000;
		Dminus[6790] = 14'b0000000_0000000;
		Dminus[6791] = 14'b0000000_0000000;
		Dminus[6792] = 14'b0000000_0000000;
		Dminus[6793] = 14'b0000000_0000000;
		Dminus[6794] = 14'b0000000_0000000;
		Dminus[6795] = 14'b0000000_0000000;
		Dminus[6796] = 14'b0000000_0000000;
		Dminus[6797] = 14'b0000000_0000000;
		Dminus[6798] = 14'b0000000_0000000;
		Dminus[6799] = 14'b0000000_0000000;
		Dminus[6800] = 14'b0000000_0000000;
		Dminus[6801] = 14'b0000000_0000000;
		Dminus[6802] = 14'b0000000_0000000;
		Dminus[6803] = 14'b0000000_0000000;
		Dminus[6804] = 14'b0000000_0000000;
		Dminus[6805] = 14'b0000000_0000000;
		Dminus[6806] = 14'b0000000_0000000;
		Dminus[6807] = 14'b0000000_0000000;
		Dminus[6808] = 14'b0000000_0000000;
		Dminus[6809] = 14'b0000000_0000000;
		Dminus[6810] = 14'b0000000_0000000;
		Dminus[6811] = 14'b0000000_0000000;
		Dminus[6812] = 14'b0000000_0000000;
		Dminus[6813] = 14'b0000000_0000000;
		Dminus[6814] = 14'b0000000_0000000;
		Dminus[6815] = 14'b0000000_0000000;
		Dminus[6816] = 14'b0000000_0000000;
		Dminus[6817] = 14'b0000000_0000000;
		Dminus[6818] = 14'b0000000_0000000;
		Dminus[6819] = 14'b0000000_0000000;
		Dminus[6820] = 14'b0000000_0000000;
		Dminus[6821] = 14'b0000000_0000000;
		Dminus[6822] = 14'b0000000_0000000;
		Dminus[6823] = 14'b0000000_0000000;
		Dminus[6824] = 14'b0000000_0000000;
		Dminus[6825] = 14'b0000000_0000000;
		Dminus[6826] = 14'b0000000_0000000;
		Dminus[6827] = 14'b0000000_0000000;
		Dminus[6828] = 14'b0000000_0000000;
		Dminus[6829] = 14'b0000000_0000000;
		Dminus[6830] = 14'b0000000_0000000;
		Dminus[6831] = 14'b0000000_0000000;
		Dminus[6832] = 14'b0000000_0000000;
		Dminus[6833] = 14'b0000000_0000000;
		Dminus[6834] = 14'b0000000_0000000;
		Dminus[6835] = 14'b0000000_0000000;
		Dminus[6836] = 14'b0000000_0000000;
		Dminus[6837] = 14'b0000000_0000000;
		Dminus[6838] = 14'b0000000_0000000;
		Dminus[6839] = 14'b0000000_0000000;
		Dminus[6840] = 14'b0000000_0000000;
		Dminus[6841] = 14'b0000000_0000000;
		Dminus[6842] = 14'b0000000_0000000;
		Dminus[6843] = 14'b0000000_0000000;
		Dminus[6844] = 14'b0000000_0000000;
		Dminus[6845] = 14'b0000000_0000000;
		Dminus[6846] = 14'b0000000_0000000;
		Dminus[6847] = 14'b0000000_0000000;
		Dminus[6848] = 14'b0000000_0000000;
		Dminus[6849] = 14'b0000000_0000000;
		Dminus[6850] = 14'b0000000_0000000;
		Dminus[6851] = 14'b0000000_0000000;
		Dminus[6852] = 14'b0000000_0000000;
		Dminus[6853] = 14'b0000000_0000000;
		Dminus[6854] = 14'b0000000_0000000;
		Dminus[6855] = 14'b0000000_0000000;
		Dminus[6856] = 14'b0000000_0000000;
		Dminus[6857] = 14'b0000000_0000000;
		Dminus[6858] = 14'b0000000_0000000;
		Dminus[6859] = 14'b0000000_0000000;
		Dminus[6860] = 14'b0000000_0000000;
		Dminus[6861] = 14'b0000000_0000000;
		Dminus[6862] = 14'b0000000_0000000;
		Dminus[6863] = 14'b0000000_0000000;
		Dminus[6864] = 14'b0000000_0000000;
		Dminus[6865] = 14'b0000000_0000000;
		Dminus[6866] = 14'b0000000_0000000;
		Dminus[6867] = 14'b0000000_0000000;
		Dminus[6868] = 14'b0000000_0000000;
		Dminus[6869] = 14'b0000000_0000000;
		Dminus[6870] = 14'b0000000_0000000;
		Dminus[6871] = 14'b0000000_0000000;
		Dminus[6872] = 14'b0000000_0000000;
		Dminus[6873] = 14'b0000000_0000000;
		Dminus[6874] = 14'b0000000_0000000;
		Dminus[6875] = 14'b0000000_0000000;
		Dminus[6876] = 14'b0000000_0000000;
		Dminus[6877] = 14'b0000000_0000000;
		Dminus[6878] = 14'b0000000_0000000;
		Dminus[6879] = 14'b0000000_0000000;
		Dminus[6880] = 14'b0000000_0000000;
		Dminus[6881] = 14'b0000000_0000000;
		Dminus[6882] = 14'b0000000_0000000;
		Dminus[6883] = 14'b0000000_0000000;
		Dminus[6884] = 14'b0000000_0000000;
		Dminus[6885] = 14'b0000000_0000000;
		Dminus[6886] = 14'b0000000_0000000;
		Dminus[6887] = 14'b0000000_0000000;
		Dminus[6888] = 14'b0000000_0000000;
		Dminus[6889] = 14'b0000000_0000000;
		Dminus[6890] = 14'b0000000_0000000;
		Dminus[6891] = 14'b0000000_0000000;
		Dminus[6892] = 14'b0000000_0000000;
		Dminus[6893] = 14'b0000000_0000000;
		Dminus[6894] = 14'b0000000_0000000;
		Dminus[6895] = 14'b0000000_0000000;
		Dminus[6896] = 14'b0000000_0000000;
		Dminus[6897] = 14'b0000000_0000000;
		Dminus[6898] = 14'b0000000_0000000;
		Dminus[6899] = 14'b0000000_0000000;
		Dminus[6900] = 14'b0000000_0000000;
		Dminus[6901] = 14'b0000000_0000000;
		Dminus[6902] = 14'b0000000_0000000;
		Dminus[6903] = 14'b0000000_0000000;
		Dminus[6904] = 14'b0000000_0000000;
		Dminus[6905] = 14'b0000000_0000000;
		Dminus[6906] = 14'b0000000_0000000;
		Dminus[6907] = 14'b0000000_0000000;
		Dminus[6908] = 14'b0000000_0000000;
		Dminus[6909] = 14'b0000000_0000000;
		Dminus[6910] = 14'b0000000_0000000;
		Dminus[6911] = 14'b0000000_0000000;
		Dminus[6912] = 14'b0000000_0000000;
		Dminus[6913] = 14'b0000000_0000000;
		Dminus[6914] = 14'b0000000_0000000;
		Dminus[6915] = 14'b0000000_0000000;
		Dminus[6916] = 14'b0000000_0000000;
		Dminus[6917] = 14'b0000000_0000000;
		Dminus[6918] = 14'b0000000_0000000;
		Dminus[6919] = 14'b0000000_0000000;
		Dminus[6920] = 14'b0000000_0000000;
		Dminus[6921] = 14'b0000000_0000000;
		Dminus[6922] = 14'b0000000_0000000;
		Dminus[6923] = 14'b0000000_0000000;
		Dminus[6924] = 14'b0000000_0000000;
		Dminus[6925] = 14'b0000000_0000000;
		Dminus[6926] = 14'b0000000_0000000;
		Dminus[6927] = 14'b0000000_0000000;
		Dminus[6928] = 14'b0000000_0000000;
		Dminus[6929] = 14'b0000000_0000000;
		Dminus[6930] = 14'b0000000_0000000;
		Dminus[6931] = 14'b0000000_0000000;
		Dminus[6932] = 14'b0000000_0000000;
		Dminus[6933] = 14'b0000000_0000000;
		Dminus[6934] = 14'b0000000_0000000;
		Dminus[6935] = 14'b0000000_0000000;
		Dminus[6936] = 14'b0000000_0000000;
		Dminus[6937] = 14'b0000000_0000000;
		Dminus[6938] = 14'b0000000_0000000;
		Dminus[6939] = 14'b0000000_0000000;
		Dminus[6940] = 14'b0000000_0000000;
		Dminus[6941] = 14'b0000000_0000000;
		Dminus[6942] = 14'b0000000_0000000;
		Dminus[6943] = 14'b0000000_0000000;
		Dminus[6944] = 14'b0000000_0000000;
		Dminus[6945] = 14'b0000000_0000000;
		Dminus[6946] = 14'b0000000_0000000;
		Dminus[6947] = 14'b0000000_0000000;
		Dminus[6948] = 14'b0000000_0000000;
		Dminus[6949] = 14'b0000000_0000000;
		Dminus[6950] = 14'b0000000_0000000;
		Dminus[6951] = 14'b0000000_0000000;
		Dminus[6952] = 14'b0000000_0000000;
		Dminus[6953] = 14'b0000000_0000000;
		Dminus[6954] = 14'b0000000_0000000;
		Dminus[6955] = 14'b0000000_0000000;
		Dminus[6956] = 14'b0000000_0000000;
		Dminus[6957] = 14'b0000000_0000000;
		Dminus[6958] = 14'b0000000_0000000;
		Dminus[6959] = 14'b0000000_0000000;
		Dminus[6960] = 14'b0000000_0000000;
		Dminus[6961] = 14'b0000000_0000000;
		Dminus[6962] = 14'b0000000_0000000;
		Dminus[6963] = 14'b0000000_0000000;
		Dminus[6964] = 14'b0000000_0000000;
		Dminus[6965] = 14'b0000000_0000000;
		Dminus[6966] = 14'b0000000_0000000;
		Dminus[6967] = 14'b0000000_0000000;
		Dminus[6968] = 14'b0000000_0000000;
		Dminus[6969] = 14'b0000000_0000000;
		Dminus[6970] = 14'b0000000_0000000;
		Dminus[6971] = 14'b0000000_0000000;
		Dminus[6972] = 14'b0000000_0000000;
		Dminus[6973] = 14'b0000000_0000000;
		Dminus[6974] = 14'b0000000_0000000;
		Dminus[6975] = 14'b0000000_0000000;
		Dminus[6976] = 14'b0000000_0000000;
		Dminus[6977] = 14'b0000000_0000000;
		Dminus[6978] = 14'b0000000_0000000;
		Dminus[6979] = 14'b0000000_0000000;
		Dminus[6980] = 14'b0000000_0000000;
		Dminus[6981] = 14'b0000000_0000000;
		Dminus[6982] = 14'b0000000_0000000;
		Dminus[6983] = 14'b0000000_0000000;
		Dminus[6984] = 14'b0000000_0000000;
		Dminus[6985] = 14'b0000000_0000000;
		Dminus[6986] = 14'b0000000_0000000;
		Dminus[6987] = 14'b0000000_0000000;
		Dminus[6988] = 14'b0000000_0000000;
		Dminus[6989] = 14'b0000000_0000000;
		Dminus[6990] = 14'b0000000_0000000;
		Dminus[6991] = 14'b0000000_0000000;
		Dminus[6992] = 14'b0000000_0000000;
		Dminus[6993] = 14'b0000000_0000000;
		Dminus[6994] = 14'b0000000_0000000;
		Dminus[6995] = 14'b0000000_0000000;
		Dminus[6996] = 14'b0000000_0000000;
		Dminus[6997] = 14'b0000000_0000000;
		Dminus[6998] = 14'b0000000_0000000;
		Dminus[6999] = 14'b0000000_0000000;
		Dminus[7000] = 14'b0000000_0000000;
		Dminus[7001] = 14'b0000000_0000000;
		Dminus[7002] = 14'b0000000_0000000;
		Dminus[7003] = 14'b0000000_0000000;
		Dminus[7004] = 14'b0000000_0000000;
		Dminus[7005] = 14'b0000000_0000000;
		Dminus[7006] = 14'b0000000_0000000;
		Dminus[7007] = 14'b0000000_0000000;
		Dminus[7008] = 14'b0000000_0000000;
		Dminus[7009] = 14'b0000000_0000000;
		Dminus[7010] = 14'b0000000_0000000;
		Dminus[7011] = 14'b0000000_0000000;
		Dminus[7012] = 14'b0000000_0000000;
		Dminus[7013] = 14'b0000000_0000000;
		Dminus[7014] = 14'b0000000_0000000;
		Dminus[7015] = 14'b0000000_0000000;
		Dminus[7016] = 14'b0000000_0000000;
		Dminus[7017] = 14'b0000000_0000000;
		Dminus[7018] = 14'b0000000_0000000;
		Dminus[7019] = 14'b0000000_0000000;
		Dminus[7020] = 14'b0000000_0000000;
		Dminus[7021] = 14'b0000000_0000000;
		Dminus[7022] = 14'b0000000_0000000;
		Dminus[7023] = 14'b0000000_0000000;
		Dminus[7024] = 14'b0000000_0000000;
		Dminus[7025] = 14'b0000000_0000000;
		Dminus[7026] = 14'b0000000_0000000;
		Dminus[7027] = 14'b0000000_0000000;
		Dminus[7028] = 14'b0000000_0000000;
		Dminus[7029] = 14'b0000000_0000000;
		Dminus[7030] = 14'b0000000_0000000;
		Dminus[7031] = 14'b0000000_0000000;
		Dminus[7032] = 14'b0000000_0000000;
		Dminus[7033] = 14'b0000000_0000000;
		Dminus[7034] = 14'b0000000_0000000;
		Dminus[7035] = 14'b0000000_0000000;
		Dminus[7036] = 14'b0000000_0000000;
		Dminus[7037] = 14'b0000000_0000000;
		Dminus[7038] = 14'b0000000_0000000;
		Dminus[7039] = 14'b0000000_0000000;
		Dminus[7040] = 14'b0000000_0000000;
		Dminus[7041] = 14'b0000000_0000000;
		Dminus[7042] = 14'b0000000_0000000;
		Dminus[7043] = 14'b0000000_0000000;
		Dminus[7044] = 14'b0000000_0000000;
		Dminus[7045] = 14'b0000000_0000000;
		Dminus[7046] = 14'b0000000_0000000;
		Dminus[7047] = 14'b0000000_0000000;
		Dminus[7048] = 14'b0000000_0000000;
		Dminus[7049] = 14'b0000000_0000000;
		Dminus[7050] = 14'b0000000_0000000;
		Dminus[7051] = 14'b0000000_0000000;
		Dminus[7052] = 14'b0000000_0000000;
		Dminus[7053] = 14'b0000000_0000000;
		Dminus[7054] = 14'b0000000_0000000;
		Dminus[7055] = 14'b0000000_0000000;
		Dminus[7056] = 14'b0000000_0000000;
		Dminus[7057] = 14'b0000000_0000000;
		Dminus[7058] = 14'b0000000_0000000;
		Dminus[7059] = 14'b0000000_0000000;
		Dminus[7060] = 14'b0000000_0000000;
		Dminus[7061] = 14'b0000000_0000000;
		Dminus[7062] = 14'b0000000_0000000;
		Dminus[7063] = 14'b0000000_0000000;
		Dminus[7064] = 14'b0000000_0000000;
		Dminus[7065] = 14'b0000000_0000000;
		Dminus[7066] = 14'b0000000_0000000;
		Dminus[7067] = 14'b0000000_0000000;
		Dminus[7068] = 14'b0000000_0000000;
		Dminus[7069] = 14'b0000000_0000000;
		Dminus[7070] = 14'b0000000_0000000;
		Dminus[7071] = 14'b0000000_0000000;
		Dminus[7072] = 14'b0000000_0000000;
		Dminus[7073] = 14'b0000000_0000000;
		Dminus[7074] = 14'b0000000_0000000;
		Dminus[7075] = 14'b0000000_0000000;
		Dminus[7076] = 14'b0000000_0000000;
		Dminus[7077] = 14'b0000000_0000000;
		Dminus[7078] = 14'b0000000_0000000;
		Dminus[7079] = 14'b0000000_0000000;
		Dminus[7080] = 14'b0000000_0000000;
		Dminus[7081] = 14'b0000000_0000000;
		Dminus[7082] = 14'b0000000_0000000;
		Dminus[7083] = 14'b0000000_0000000;
		Dminus[7084] = 14'b0000000_0000000;
		Dminus[7085] = 14'b0000000_0000000;
		Dminus[7086] = 14'b0000000_0000000;
		Dminus[7087] = 14'b0000000_0000000;
		Dminus[7088] = 14'b0000000_0000000;
		Dminus[7089] = 14'b0000000_0000000;
		Dminus[7090] = 14'b0000000_0000000;
		Dminus[7091] = 14'b0000000_0000000;
		Dminus[7092] = 14'b0000000_0000000;
		Dminus[7093] = 14'b0000000_0000000;
		Dminus[7094] = 14'b0000000_0000000;
		Dminus[7095] = 14'b0000000_0000000;
		Dminus[7096] = 14'b0000000_0000000;
		Dminus[7097] = 14'b0000000_0000000;
		Dminus[7098] = 14'b0000000_0000000;
		Dminus[7099] = 14'b0000000_0000000;
		Dminus[7100] = 14'b0000000_0000000;
		Dminus[7101] = 14'b0000000_0000000;
		Dminus[7102] = 14'b0000000_0000000;
		Dminus[7103] = 14'b0000000_0000000;
		Dminus[7104] = 14'b0000000_0000000;
		Dminus[7105] = 14'b0000000_0000000;
		Dminus[7106] = 14'b0000000_0000000;
		Dminus[7107] = 14'b0000000_0000000;
		Dminus[7108] = 14'b0000000_0000000;
		Dminus[7109] = 14'b0000000_0000000;
		Dminus[7110] = 14'b0000000_0000000;
		Dminus[7111] = 14'b0000000_0000000;
		Dminus[7112] = 14'b0000000_0000000;
		Dminus[7113] = 14'b0000000_0000000;
		Dminus[7114] = 14'b0000000_0000000;
		Dminus[7115] = 14'b0000000_0000000;
		Dminus[7116] = 14'b0000000_0000000;
		Dminus[7117] = 14'b0000000_0000000;
		Dminus[7118] = 14'b0000000_0000000;
		Dminus[7119] = 14'b0000000_0000000;
		Dminus[7120] = 14'b0000000_0000000;
		Dminus[7121] = 14'b0000000_0000000;
		Dminus[7122] = 14'b0000000_0000000;
		Dminus[7123] = 14'b0000000_0000000;
		Dminus[7124] = 14'b0000000_0000000;
		Dminus[7125] = 14'b0000000_0000000;
		Dminus[7126] = 14'b0000000_0000000;
		Dminus[7127] = 14'b0000000_0000000;
		Dminus[7128] = 14'b0000000_0000000;
		Dminus[7129] = 14'b0000000_0000000;
		Dminus[7130] = 14'b0000000_0000000;
		Dminus[7131] = 14'b0000000_0000000;
		Dminus[7132] = 14'b0000000_0000000;
		Dminus[7133] = 14'b0000000_0000000;
		Dminus[7134] = 14'b0000000_0000000;
		Dminus[7135] = 14'b0000000_0000000;
		Dminus[7136] = 14'b0000000_0000000;
		Dminus[7137] = 14'b0000000_0000000;
		Dminus[7138] = 14'b0000000_0000000;
		Dminus[7139] = 14'b0000000_0000000;
		Dminus[7140] = 14'b0000000_0000000;
		Dminus[7141] = 14'b0000000_0000000;
		Dminus[7142] = 14'b0000000_0000000;
		Dminus[7143] = 14'b0000000_0000000;
		Dminus[7144] = 14'b0000000_0000000;
		Dminus[7145] = 14'b0000000_0000000;
		Dminus[7146] = 14'b0000000_0000000;
		Dminus[7147] = 14'b0000000_0000000;
		Dminus[7148] = 14'b0000000_0000000;
		Dminus[7149] = 14'b0000000_0000000;
		Dminus[7150] = 14'b0000000_0000000;
		Dminus[7151] = 14'b0000000_0000000;
		Dminus[7152] = 14'b0000000_0000000;
		Dminus[7153] = 14'b0000000_0000000;
		Dminus[7154] = 14'b0000000_0000000;
		Dminus[7155] = 14'b0000000_0000000;
		Dminus[7156] = 14'b0000000_0000000;
		Dminus[7157] = 14'b0000000_0000000;
		Dminus[7158] = 14'b0000000_0000000;
		Dminus[7159] = 14'b0000000_0000000;
		Dminus[7160] = 14'b0000000_0000000;
		Dminus[7161] = 14'b0000000_0000000;
		Dminus[7162] = 14'b0000000_0000000;
		Dminus[7163] = 14'b0000000_0000000;
		Dminus[7164] = 14'b0000000_0000000;
		Dminus[7165] = 14'b0000000_0000000;
		Dminus[7166] = 14'b0000000_0000000;
		Dminus[7167] = 14'b0000000_0000000;
		Dminus[7168] = 14'b0000000_0000000;
		Dminus[7169] = 14'b0000000_0000000;
		Dminus[7170] = 14'b0000000_0000000;
		Dminus[7171] = 14'b0000000_0000000;
		Dminus[7172] = 14'b0000000_0000000;
		Dminus[7173] = 14'b0000000_0000000;
		Dminus[7174] = 14'b0000000_0000000;
		Dminus[7175] = 14'b0000000_0000000;
		Dminus[7176] = 14'b0000000_0000000;
		Dminus[7177] = 14'b0000000_0000000;
		Dminus[7178] = 14'b0000000_0000000;
		Dminus[7179] = 14'b0000000_0000000;
		Dminus[7180] = 14'b0000000_0000000;
		Dminus[7181] = 14'b0000000_0000000;
		Dminus[7182] = 14'b0000000_0000000;
		Dminus[7183] = 14'b0000000_0000000;
		Dminus[7184] = 14'b0000000_0000000;
		Dminus[7185] = 14'b0000000_0000000;
		Dminus[7186] = 14'b0000000_0000000;
		Dminus[7187] = 14'b0000000_0000000;
		Dminus[7188] = 14'b0000000_0000000;
		Dminus[7189] = 14'b0000000_0000000;
		Dminus[7190] = 14'b0000000_0000000;
		Dminus[7191] = 14'b0000000_0000000;
		Dminus[7192] = 14'b0000000_0000000;
		Dminus[7193] = 14'b0000000_0000000;
		Dminus[7194] = 14'b0000000_0000000;
		Dminus[7195] = 14'b0000000_0000000;
		Dminus[7196] = 14'b0000000_0000000;
		Dminus[7197] = 14'b0000000_0000000;
		Dminus[7198] = 14'b0000000_0000000;
		Dminus[7199] = 14'b0000000_0000000;
		Dminus[7200] = 14'b0000000_0000000;
		Dminus[7201] = 14'b0000000_0000000;
		Dminus[7202] = 14'b0000000_0000000;
		Dminus[7203] = 14'b0000000_0000000;
		Dminus[7204] = 14'b0000000_0000000;
		Dminus[7205] = 14'b0000000_0000000;
		Dminus[7206] = 14'b0000000_0000000;
		Dminus[7207] = 14'b0000000_0000000;
		Dminus[7208] = 14'b0000000_0000000;
		Dminus[7209] = 14'b0000000_0000000;
		Dminus[7210] = 14'b0000000_0000000;
		Dminus[7211] = 14'b0000000_0000000;
		Dminus[7212] = 14'b0000000_0000000;
		Dminus[7213] = 14'b0000000_0000000;
		Dminus[7214] = 14'b0000000_0000000;
		Dminus[7215] = 14'b0000000_0000000;
		Dminus[7216] = 14'b0000000_0000000;
		Dminus[7217] = 14'b0000000_0000000;
		Dminus[7218] = 14'b0000000_0000000;
		Dminus[7219] = 14'b0000000_0000000;
		Dminus[7220] = 14'b0000000_0000000;
		Dminus[7221] = 14'b0000000_0000000;
		Dminus[7222] = 14'b0000000_0000000;
		Dminus[7223] = 14'b0000000_0000000;
		Dminus[7224] = 14'b0000000_0000000;
		Dminus[7225] = 14'b0000000_0000000;
		Dminus[7226] = 14'b0000000_0000000;
		Dminus[7227] = 14'b0000000_0000000;
		Dminus[7228] = 14'b0000000_0000000;
		Dminus[7229] = 14'b0000000_0000000;
		Dminus[7230] = 14'b0000000_0000000;
		Dminus[7231] = 14'b0000000_0000000;
		Dminus[7232] = 14'b0000000_0000000;
		Dminus[7233] = 14'b0000000_0000000;
		Dminus[7234] = 14'b0000000_0000000;
		Dminus[7235] = 14'b0000000_0000000;
		Dminus[7236] = 14'b0000000_0000000;
		Dminus[7237] = 14'b0000000_0000000;
		Dminus[7238] = 14'b0000000_0000000;
		Dminus[7239] = 14'b0000000_0000000;
		Dminus[7240] = 14'b0000000_0000000;
		Dminus[7241] = 14'b0000000_0000000;
		Dminus[7242] = 14'b0000000_0000000;
		Dminus[7243] = 14'b0000000_0000000;
		Dminus[7244] = 14'b0000000_0000000;
		Dminus[7245] = 14'b0000000_0000000;
		Dminus[7246] = 14'b0000000_0000000;
		Dminus[7247] = 14'b0000000_0000000;
		Dminus[7248] = 14'b0000000_0000000;
		Dminus[7249] = 14'b0000000_0000000;
		Dminus[7250] = 14'b0000000_0000000;
		Dminus[7251] = 14'b0000000_0000000;
		Dminus[7252] = 14'b0000000_0000000;
		Dminus[7253] = 14'b0000000_0000000;
		Dminus[7254] = 14'b0000000_0000000;
		Dminus[7255] = 14'b0000000_0000000;
		Dminus[7256] = 14'b0000000_0000000;
		Dminus[7257] = 14'b0000000_0000000;
		Dminus[7258] = 14'b0000000_0000000;
		Dminus[7259] = 14'b0000000_0000000;
		Dminus[7260] = 14'b0000000_0000000;
		Dminus[7261] = 14'b0000000_0000000;
		Dminus[7262] = 14'b0000000_0000000;
		Dminus[7263] = 14'b0000000_0000000;
		Dminus[7264] = 14'b0000000_0000000;
		Dminus[7265] = 14'b0000000_0000000;
		Dminus[7266] = 14'b0000000_0000000;
		Dminus[7267] = 14'b0000000_0000000;
		Dminus[7268] = 14'b0000000_0000000;
		Dminus[7269] = 14'b0000000_0000000;
		Dminus[7270] = 14'b0000000_0000000;
		Dminus[7271] = 14'b0000000_0000000;
		Dminus[7272] = 14'b0000000_0000000;
		Dminus[7273] = 14'b0000000_0000000;
		Dminus[7274] = 14'b0000000_0000000;
		Dminus[7275] = 14'b0000000_0000000;
		Dminus[7276] = 14'b0000000_0000000;
		Dminus[7277] = 14'b0000000_0000000;
		Dminus[7278] = 14'b0000000_0000000;
		Dminus[7279] = 14'b0000000_0000000;
		Dminus[7280] = 14'b0000000_0000000;
		Dminus[7281] = 14'b0000000_0000000;
		Dminus[7282] = 14'b0000000_0000000;
		Dminus[7283] = 14'b0000000_0000000;
		Dminus[7284] = 14'b0000000_0000000;
		Dminus[7285] = 14'b0000000_0000000;
		Dminus[7286] = 14'b0000000_0000000;
		Dminus[7287] = 14'b0000000_0000000;
		Dminus[7288] = 14'b0000000_0000000;
		Dminus[7289] = 14'b0000000_0000000;
		Dminus[7290] = 14'b0000000_0000000;
		Dminus[7291] = 14'b0000000_0000000;
		Dminus[7292] = 14'b0000000_0000000;
		Dminus[7293] = 14'b0000000_0000000;
		Dminus[7294] = 14'b0000000_0000000;
		Dminus[7295] = 14'b0000000_0000000;
		Dminus[7296] = 14'b0000000_0000000;
		Dminus[7297] = 14'b0000000_0000000;
		Dminus[7298] = 14'b0000000_0000000;
		Dminus[7299] = 14'b0000000_0000000;
		Dminus[7300] = 14'b0000000_0000000;
		Dminus[7301] = 14'b0000000_0000000;
		Dminus[7302] = 14'b0000000_0000000;
		Dminus[7303] = 14'b0000000_0000000;
		Dminus[7304] = 14'b0000000_0000000;
		Dminus[7305] = 14'b0000000_0000000;
		Dminus[7306] = 14'b0000000_0000000;
		Dminus[7307] = 14'b0000000_0000000;
		Dminus[7308] = 14'b0000000_0000000;
		Dminus[7309] = 14'b0000000_0000000;
		Dminus[7310] = 14'b0000000_0000000;
		Dminus[7311] = 14'b0000000_0000000;
		Dminus[7312] = 14'b0000000_0000000;
		Dminus[7313] = 14'b0000000_0000000;
		Dminus[7314] = 14'b0000000_0000000;
		Dminus[7315] = 14'b0000000_0000000;
		Dminus[7316] = 14'b0000000_0000000;
		Dminus[7317] = 14'b0000000_0000000;
		Dminus[7318] = 14'b0000000_0000000;
		Dminus[7319] = 14'b0000000_0000000;
		Dminus[7320] = 14'b0000000_0000000;
		Dminus[7321] = 14'b0000000_0000000;
		Dminus[7322] = 14'b0000000_0000000;
		Dminus[7323] = 14'b0000000_0000000;
		Dminus[7324] = 14'b0000000_0000000;
		Dminus[7325] = 14'b0000000_0000000;
		Dminus[7326] = 14'b0000000_0000000;
		Dminus[7327] = 14'b0000000_0000000;
		Dminus[7328] = 14'b0000000_0000000;
		Dminus[7329] = 14'b0000000_0000000;
		Dminus[7330] = 14'b0000000_0000000;
		Dminus[7331] = 14'b0000000_0000000;
		Dminus[7332] = 14'b0000000_0000000;
		Dminus[7333] = 14'b0000000_0000000;
		Dminus[7334] = 14'b0000000_0000000;
		Dminus[7335] = 14'b0000000_0000000;
		Dminus[7336] = 14'b0000000_0000000;
		Dminus[7337] = 14'b0000000_0000000;
		Dminus[7338] = 14'b0000000_0000000;
		Dminus[7339] = 14'b0000000_0000000;
		Dminus[7340] = 14'b0000000_0000000;
		Dminus[7341] = 14'b0000000_0000000;
		Dminus[7342] = 14'b0000000_0000000;
		Dminus[7343] = 14'b0000000_0000000;
		Dminus[7344] = 14'b0000000_0000000;
		Dminus[7345] = 14'b0000000_0000000;
		Dminus[7346] = 14'b0000000_0000000;
		Dminus[7347] = 14'b0000000_0000000;
		Dminus[7348] = 14'b0000000_0000000;
		Dminus[7349] = 14'b0000000_0000000;
		Dminus[7350] = 14'b0000000_0000000;
		Dminus[7351] = 14'b0000000_0000000;
		Dminus[7352] = 14'b0000000_0000000;
		Dminus[7353] = 14'b0000000_0000000;
		Dminus[7354] = 14'b0000000_0000000;
		Dminus[7355] = 14'b0000000_0000000;
		Dminus[7356] = 14'b0000000_0000000;
		Dminus[7357] = 14'b0000000_0000000;
		Dminus[7358] = 14'b0000000_0000000;
		Dminus[7359] = 14'b0000000_0000000;
		Dminus[7360] = 14'b0000000_0000000;
		Dminus[7361] = 14'b0000000_0000000;
		Dminus[7362] = 14'b0000000_0000000;
		Dminus[7363] = 14'b0000000_0000000;
		Dminus[7364] = 14'b0000000_0000000;
		Dminus[7365] = 14'b0000000_0000000;
		Dminus[7366] = 14'b0000000_0000000;
		Dminus[7367] = 14'b0000000_0000000;
		Dminus[7368] = 14'b0000000_0000000;
		Dminus[7369] = 14'b0000000_0000000;
		Dminus[7370] = 14'b0000000_0000000;
		Dminus[7371] = 14'b0000000_0000000;
		Dminus[7372] = 14'b0000000_0000000;
		Dminus[7373] = 14'b0000000_0000000;
		Dminus[7374] = 14'b0000000_0000000;
		Dminus[7375] = 14'b0000000_0000000;
		Dminus[7376] = 14'b0000000_0000000;
		Dminus[7377] = 14'b0000000_0000000;
		Dminus[7378] = 14'b0000000_0000000;
		Dminus[7379] = 14'b0000000_0000000;
		Dminus[7380] = 14'b0000000_0000000;
		Dminus[7381] = 14'b0000000_0000000;
		Dminus[7382] = 14'b0000000_0000000;
		Dminus[7383] = 14'b0000000_0000000;
		Dminus[7384] = 14'b0000000_0000000;
		Dminus[7385] = 14'b0000000_0000000;
		Dminus[7386] = 14'b0000000_0000000;
		Dminus[7387] = 14'b0000000_0000000;
		Dminus[7388] = 14'b0000000_0000000;
		Dminus[7389] = 14'b0000000_0000000;
		Dminus[7390] = 14'b0000000_0000000;
		Dminus[7391] = 14'b0000000_0000000;
		Dminus[7392] = 14'b0000000_0000000;
		Dminus[7393] = 14'b0000000_0000000;
		Dminus[7394] = 14'b0000000_0000000;
		Dminus[7395] = 14'b0000000_0000000;
		Dminus[7396] = 14'b0000000_0000000;
		Dminus[7397] = 14'b0000000_0000000;
		Dminus[7398] = 14'b0000000_0000000;
		Dminus[7399] = 14'b0000000_0000000;
		Dminus[7400] = 14'b0000000_0000000;
		Dminus[7401] = 14'b0000000_0000000;
		Dminus[7402] = 14'b0000000_0000000;
		Dminus[7403] = 14'b0000000_0000000;
		Dminus[7404] = 14'b0000000_0000000;
		Dminus[7405] = 14'b0000000_0000000;
		Dminus[7406] = 14'b0000000_0000000;
		Dminus[7407] = 14'b0000000_0000000;
		Dminus[7408] = 14'b0000000_0000000;
		Dminus[7409] = 14'b0000000_0000000;
		Dminus[7410] = 14'b0000000_0000000;
		Dminus[7411] = 14'b0000000_0000000;
		Dminus[7412] = 14'b0000000_0000000;
		Dminus[7413] = 14'b0000000_0000000;
		Dminus[7414] = 14'b0000000_0000000;
		Dminus[7415] = 14'b0000000_0000000;
		Dminus[7416] = 14'b0000000_0000000;
		Dminus[7417] = 14'b0000000_0000000;
		Dminus[7418] = 14'b0000000_0000000;
		Dminus[7419] = 14'b0000000_0000000;
		Dminus[7420] = 14'b0000000_0000000;
		Dminus[7421] = 14'b0000000_0000000;
		Dminus[7422] = 14'b0000000_0000000;
		Dminus[7423] = 14'b0000000_0000000;
		Dminus[7424] = 14'b0000000_0000000;
		Dminus[7425] = 14'b0000000_0000000;
		Dminus[7426] = 14'b0000000_0000000;
		Dminus[7427] = 14'b0000000_0000000;
		Dminus[7428] = 14'b0000000_0000000;
		Dminus[7429] = 14'b0000000_0000000;
		Dminus[7430] = 14'b0000000_0000000;
		Dminus[7431] = 14'b0000000_0000000;
		Dminus[7432] = 14'b0000000_0000000;
		Dminus[7433] = 14'b0000000_0000000;
		Dminus[7434] = 14'b0000000_0000000;
		Dminus[7435] = 14'b0000000_0000000;
		Dminus[7436] = 14'b0000000_0000000;
		Dminus[7437] = 14'b0000000_0000000;
		Dminus[7438] = 14'b0000000_0000000;
		Dminus[7439] = 14'b0000000_0000000;
		Dminus[7440] = 14'b0000000_0000000;
		Dminus[7441] = 14'b0000000_0000000;
		Dminus[7442] = 14'b0000000_0000000;
		Dminus[7443] = 14'b0000000_0000000;
		Dminus[7444] = 14'b0000000_0000000;
		Dminus[7445] = 14'b0000000_0000000;
		Dminus[7446] = 14'b0000000_0000000;
		Dminus[7447] = 14'b0000000_0000000;
		Dminus[7448] = 14'b0000000_0000000;
		Dminus[7449] = 14'b0000000_0000000;
		Dminus[7450] = 14'b0000000_0000000;
		Dminus[7451] = 14'b0000000_0000000;
		Dminus[7452] = 14'b0000000_0000000;
		Dminus[7453] = 14'b0000000_0000000;
		Dminus[7454] = 14'b0000000_0000000;
		Dminus[7455] = 14'b0000000_0000000;
		Dminus[7456] = 14'b0000000_0000000;
		Dminus[7457] = 14'b0000000_0000000;
		Dminus[7458] = 14'b0000000_0000000;
		Dminus[7459] = 14'b0000000_0000000;
		Dminus[7460] = 14'b0000000_0000000;
		Dminus[7461] = 14'b0000000_0000000;
		Dminus[7462] = 14'b0000000_0000000;
		Dminus[7463] = 14'b0000000_0000000;
		Dminus[7464] = 14'b0000000_0000000;
		Dminus[7465] = 14'b0000000_0000000;
		Dminus[7466] = 14'b0000000_0000000;
		Dminus[7467] = 14'b0000000_0000000;
		Dminus[7468] = 14'b0000000_0000000;
		Dminus[7469] = 14'b0000000_0000000;
		Dminus[7470] = 14'b0000000_0000000;
		Dminus[7471] = 14'b0000000_0000000;
		Dminus[7472] = 14'b0000000_0000000;
		Dminus[7473] = 14'b0000000_0000000;
		Dminus[7474] = 14'b0000000_0000000;
		Dminus[7475] = 14'b0000000_0000000;
		Dminus[7476] = 14'b0000000_0000000;
		Dminus[7477] = 14'b0000000_0000000;
		Dminus[7478] = 14'b0000000_0000000;
		Dminus[7479] = 14'b0000000_0000000;
		Dminus[7480] = 14'b0000000_0000000;
		Dminus[7481] = 14'b0000000_0000000;
		Dminus[7482] = 14'b0000000_0000000;
		Dminus[7483] = 14'b0000000_0000000;
		Dminus[7484] = 14'b0000000_0000000;
		Dminus[7485] = 14'b0000000_0000000;
		Dminus[7486] = 14'b0000000_0000000;
		Dminus[7487] = 14'b0000000_0000000;
		Dminus[7488] = 14'b0000000_0000000;
		Dminus[7489] = 14'b0000000_0000000;
		Dminus[7490] = 14'b0000000_0000000;
		Dminus[7491] = 14'b0000000_0000000;
		Dminus[7492] = 14'b0000000_0000000;
		Dminus[7493] = 14'b0000000_0000000;
		Dminus[7494] = 14'b0000000_0000000;
		Dminus[7495] = 14'b0000000_0000000;
		Dminus[7496] = 14'b0000000_0000000;
		Dminus[7497] = 14'b0000000_0000000;
		Dminus[7498] = 14'b0000000_0000000;
		Dminus[7499] = 14'b0000000_0000000;
		Dminus[7500] = 14'b0000000_0000000;
		Dminus[7501] = 14'b0000000_0000000;
		Dminus[7502] = 14'b0000000_0000000;
		Dminus[7503] = 14'b0000000_0000000;
		Dminus[7504] = 14'b0000000_0000000;
		Dminus[7505] = 14'b0000000_0000000;
		Dminus[7506] = 14'b0000000_0000000;
		Dminus[7507] = 14'b0000000_0000000;
		Dminus[7508] = 14'b0000000_0000000;
		Dminus[7509] = 14'b0000000_0000000;
		Dminus[7510] = 14'b0000000_0000000;
		Dminus[7511] = 14'b0000000_0000000;
		Dminus[7512] = 14'b0000000_0000000;
		Dminus[7513] = 14'b0000000_0000000;
		Dminus[7514] = 14'b0000000_0000000;
		Dminus[7515] = 14'b0000000_0000000;
		Dminus[7516] = 14'b0000000_0000000;
		Dminus[7517] = 14'b0000000_0000000;
		Dminus[7518] = 14'b0000000_0000000;
		Dminus[7519] = 14'b0000000_0000000;
		Dminus[7520] = 14'b0000000_0000000;
		Dminus[7521] = 14'b0000000_0000000;
		Dminus[7522] = 14'b0000000_0000000;
		Dminus[7523] = 14'b0000000_0000000;
		Dminus[7524] = 14'b0000000_0000000;
		Dminus[7525] = 14'b0000000_0000000;
		Dminus[7526] = 14'b0000000_0000000;
		Dminus[7527] = 14'b0000000_0000000;
		Dminus[7528] = 14'b0000000_0000000;
		Dminus[7529] = 14'b0000000_0000000;
		Dminus[7530] = 14'b0000000_0000000;
		Dminus[7531] = 14'b0000000_0000000;
		Dminus[7532] = 14'b0000000_0000000;
		Dminus[7533] = 14'b0000000_0000000;
		Dminus[7534] = 14'b0000000_0000000;
		Dminus[7535] = 14'b0000000_0000000;
		Dminus[7536] = 14'b0000000_0000000;
		Dminus[7537] = 14'b0000000_0000000;
		Dminus[7538] = 14'b0000000_0000000;
		Dminus[7539] = 14'b0000000_0000000;
		Dminus[7540] = 14'b0000000_0000000;
		Dminus[7541] = 14'b0000000_0000000;
		Dminus[7542] = 14'b0000000_0000000;
		Dminus[7543] = 14'b0000000_0000000;
		Dminus[7544] = 14'b0000000_0000000;
		Dminus[7545] = 14'b0000000_0000000;
		Dminus[7546] = 14'b0000000_0000000;
		Dminus[7547] = 14'b0000000_0000000;
		Dminus[7548] = 14'b0000000_0000000;
		Dminus[7549] = 14'b0000000_0000000;
		Dminus[7550] = 14'b0000000_0000000;
		Dminus[7551] = 14'b0000000_0000000;
		Dminus[7552] = 14'b0000000_0000000;
		Dminus[7553] = 14'b0000000_0000000;
		Dminus[7554] = 14'b0000000_0000000;
		Dminus[7555] = 14'b0000000_0000000;
		Dminus[7556] = 14'b0000000_0000000;
		Dminus[7557] = 14'b0000000_0000000;
		Dminus[7558] = 14'b0000000_0000000;
		Dminus[7559] = 14'b0000000_0000000;
		Dminus[7560] = 14'b0000000_0000000;
		Dminus[7561] = 14'b0000000_0000000;
		Dminus[7562] = 14'b0000000_0000000;
		Dminus[7563] = 14'b0000000_0000000;
		Dminus[7564] = 14'b0000000_0000000;
		Dminus[7565] = 14'b0000000_0000000;
		Dminus[7566] = 14'b0000000_0000000;
		Dminus[7567] = 14'b0000000_0000000;
		Dminus[7568] = 14'b0000000_0000000;
		Dminus[7569] = 14'b0000000_0000000;
		Dminus[7570] = 14'b0000000_0000000;
		Dminus[7571] = 14'b0000000_0000000;
		Dminus[7572] = 14'b0000000_0000000;
		Dminus[7573] = 14'b0000000_0000000;
		Dminus[7574] = 14'b0000000_0000000;
		Dminus[7575] = 14'b0000000_0000000;
		Dminus[7576] = 14'b0000000_0000000;
		Dminus[7577] = 14'b0000000_0000000;
		Dminus[7578] = 14'b0000000_0000000;
		Dminus[7579] = 14'b0000000_0000000;
		Dminus[7580] = 14'b0000000_0000000;
		Dminus[7581] = 14'b0000000_0000000;
		Dminus[7582] = 14'b0000000_0000000;
		Dminus[7583] = 14'b0000000_0000000;
		Dminus[7584] = 14'b0000000_0000000;
		Dminus[7585] = 14'b0000000_0000000;
		Dminus[7586] = 14'b0000000_0000000;
		Dminus[7587] = 14'b0000000_0000000;
		Dminus[7588] = 14'b0000000_0000000;
		Dminus[7589] = 14'b0000000_0000000;
		Dminus[7590] = 14'b0000000_0000000;
		Dminus[7591] = 14'b0000000_0000000;
		Dminus[7592] = 14'b0000000_0000000;
		Dminus[7593] = 14'b0000000_0000000;
		Dminus[7594] = 14'b0000000_0000000;
		Dminus[7595] = 14'b0000000_0000000;
		Dminus[7596] = 14'b0000000_0000000;
		Dminus[7597] = 14'b0000000_0000000;
		Dminus[7598] = 14'b0000000_0000000;
		Dminus[7599] = 14'b0000000_0000000;
		Dminus[7600] = 14'b0000000_0000000;
		Dminus[7601] = 14'b0000000_0000000;
		Dminus[7602] = 14'b0000000_0000000;
		Dminus[7603] = 14'b0000000_0000000;
		Dminus[7604] = 14'b0000000_0000000;
		Dminus[7605] = 14'b0000000_0000000;
		Dminus[7606] = 14'b0000000_0000000;
		Dminus[7607] = 14'b0000000_0000000;
		Dminus[7608] = 14'b0000000_0000000;
		Dminus[7609] = 14'b0000000_0000000;
		Dminus[7610] = 14'b0000000_0000000;
		Dminus[7611] = 14'b0000000_0000000;
		Dminus[7612] = 14'b0000000_0000000;
		Dminus[7613] = 14'b0000000_0000000;
		Dminus[7614] = 14'b0000000_0000000;
		Dminus[7615] = 14'b0000000_0000000;
		Dminus[7616] = 14'b0000000_0000000;
		Dminus[7617] = 14'b0000000_0000000;
		Dminus[7618] = 14'b0000000_0000000;
		Dminus[7619] = 14'b0000000_0000000;
		Dminus[7620] = 14'b0000000_0000000;
		Dminus[7621] = 14'b0000000_0000000;
		Dminus[7622] = 14'b0000000_0000000;
		Dminus[7623] = 14'b0000000_0000000;
		Dminus[7624] = 14'b0000000_0000000;
		Dminus[7625] = 14'b0000000_0000000;
		Dminus[7626] = 14'b0000000_0000000;
		Dminus[7627] = 14'b0000000_0000000;
		Dminus[7628] = 14'b0000000_0000000;
		Dminus[7629] = 14'b0000000_0000000;
		Dminus[7630] = 14'b0000000_0000000;
		Dminus[7631] = 14'b0000000_0000000;
		Dminus[7632] = 14'b0000000_0000000;
		Dminus[7633] = 14'b0000000_0000000;
		Dminus[7634] = 14'b0000000_0000000;
		Dminus[7635] = 14'b0000000_0000000;
		Dminus[7636] = 14'b0000000_0000000;
		Dminus[7637] = 14'b0000000_0000000;
		Dminus[7638] = 14'b0000000_0000000;
		Dminus[7639] = 14'b0000000_0000000;
		Dminus[7640] = 14'b0000000_0000000;
		Dminus[7641] = 14'b0000000_0000000;
		Dminus[7642] = 14'b0000000_0000000;
		Dminus[7643] = 14'b0000000_0000000;
		Dminus[7644] = 14'b0000000_0000000;
		Dminus[7645] = 14'b0000000_0000000;
		Dminus[7646] = 14'b0000000_0000000;
		Dminus[7647] = 14'b0000000_0000000;
		Dminus[7648] = 14'b0000000_0000000;
		Dminus[7649] = 14'b0000000_0000000;
		Dminus[7650] = 14'b0000000_0000000;
		Dminus[7651] = 14'b0000000_0000000;
		Dminus[7652] = 14'b0000000_0000000;
		Dminus[7653] = 14'b0000000_0000000;
		Dminus[7654] = 14'b0000000_0000000;
		Dminus[7655] = 14'b0000000_0000000;
		Dminus[7656] = 14'b0000000_0000000;
		Dminus[7657] = 14'b0000000_0000000;
		Dminus[7658] = 14'b0000000_0000000;
		Dminus[7659] = 14'b0000000_0000000;
		Dminus[7660] = 14'b0000000_0000000;
		Dminus[7661] = 14'b0000000_0000000;
		Dminus[7662] = 14'b0000000_0000000;
		Dminus[7663] = 14'b0000000_0000000;
		Dminus[7664] = 14'b0000000_0000000;
		Dminus[7665] = 14'b0000000_0000000;
		Dminus[7666] = 14'b0000000_0000000;
		Dminus[7667] = 14'b0000000_0000000;
		Dminus[7668] = 14'b0000000_0000000;
		Dminus[7669] = 14'b0000000_0000000;
		Dminus[7670] = 14'b0000000_0000000;
		Dminus[7671] = 14'b0000000_0000000;
		Dminus[7672] = 14'b0000000_0000000;
		Dminus[7673] = 14'b0000000_0000000;
		Dminus[7674] = 14'b0000000_0000000;
		Dminus[7675] = 14'b0000000_0000000;
		Dminus[7676] = 14'b0000000_0000000;
		Dminus[7677] = 14'b0000000_0000000;
		Dminus[7678] = 14'b0000000_0000000;
		Dminus[7679] = 14'b0000000_0000000;
		Dminus[7680] = 14'b0000000_0000000;
		Dminus[7681] = 14'b0000000_0000000;
		Dminus[7682] = 14'b0000000_0000000;
		Dminus[7683] = 14'b0000000_0000000;
		Dminus[7684] = 14'b0000000_0000000;
		Dminus[7685] = 14'b0000000_0000000;
		Dminus[7686] = 14'b0000000_0000000;
		Dminus[7687] = 14'b0000000_0000000;
		Dminus[7688] = 14'b0000000_0000000;
		Dminus[7689] = 14'b0000000_0000000;
		Dminus[7690] = 14'b0000000_0000000;
		Dminus[7691] = 14'b0000000_0000000;
		Dminus[7692] = 14'b0000000_0000000;
		Dminus[7693] = 14'b0000000_0000000;
		Dminus[7694] = 14'b0000000_0000000;
		Dminus[7695] = 14'b0000000_0000000;
		Dminus[7696] = 14'b0000000_0000000;
		Dminus[7697] = 14'b0000000_0000000;
		Dminus[7698] = 14'b0000000_0000000;
		Dminus[7699] = 14'b0000000_0000000;
		Dminus[7700] = 14'b0000000_0000000;
		Dminus[7701] = 14'b0000000_0000000;
		Dminus[7702] = 14'b0000000_0000000;
		Dminus[7703] = 14'b0000000_0000000;
		Dminus[7704] = 14'b0000000_0000000;
		Dminus[7705] = 14'b0000000_0000000;
		Dminus[7706] = 14'b0000000_0000000;
		Dminus[7707] = 14'b0000000_0000000;
		Dminus[7708] = 14'b0000000_0000000;
		Dminus[7709] = 14'b0000000_0000000;
		Dminus[7710] = 14'b0000000_0000000;
		Dminus[7711] = 14'b0000000_0000000;
		Dminus[7712] = 14'b0000000_0000000;
		Dminus[7713] = 14'b0000000_0000000;
		Dminus[7714] = 14'b0000000_0000000;
		Dminus[7715] = 14'b0000000_0000000;
		Dminus[7716] = 14'b0000000_0000000;
		Dminus[7717] = 14'b0000000_0000000;
		Dminus[7718] = 14'b0000000_0000000;
		Dminus[7719] = 14'b0000000_0000000;
		Dminus[7720] = 14'b0000000_0000000;
		Dminus[7721] = 14'b0000000_0000000;
		Dminus[7722] = 14'b0000000_0000000;
		Dminus[7723] = 14'b0000000_0000000;
		Dminus[7724] = 14'b0000000_0000000;
		Dminus[7725] = 14'b0000000_0000000;
		Dminus[7726] = 14'b0000000_0000000;
		Dminus[7727] = 14'b0000000_0000000;
		Dminus[7728] = 14'b0000000_0000000;
		Dminus[7729] = 14'b0000000_0000000;
		Dminus[7730] = 14'b0000000_0000000;
		Dminus[7731] = 14'b0000000_0000000;
		Dminus[7732] = 14'b0000000_0000000;
		Dminus[7733] = 14'b0000000_0000000;
		Dminus[7734] = 14'b0000000_0000000;
		Dminus[7735] = 14'b0000000_0000000;
		Dminus[7736] = 14'b0000000_0000000;
		Dminus[7737] = 14'b0000000_0000000;
		Dminus[7738] = 14'b0000000_0000000;
		Dminus[7739] = 14'b0000000_0000000;
		Dminus[7740] = 14'b0000000_0000000;
		Dminus[7741] = 14'b0000000_0000000;
		Dminus[7742] = 14'b0000000_0000000;
		Dminus[7743] = 14'b0000000_0000000;
		Dminus[7744] = 14'b0000000_0000000;
		Dminus[7745] = 14'b0000000_0000000;
		Dminus[7746] = 14'b0000000_0000000;
		Dminus[7747] = 14'b0000000_0000000;
		Dminus[7748] = 14'b0000000_0000000;
		Dminus[7749] = 14'b0000000_0000000;
		Dminus[7750] = 14'b0000000_0000000;
		Dminus[7751] = 14'b0000000_0000000;
		Dminus[7752] = 14'b0000000_0000000;
		Dminus[7753] = 14'b0000000_0000000;
		Dminus[7754] = 14'b0000000_0000000;
		Dminus[7755] = 14'b0000000_0000000;
		Dminus[7756] = 14'b0000000_0000000;
		Dminus[7757] = 14'b0000000_0000000;
		Dminus[7758] = 14'b0000000_0000000;
		Dminus[7759] = 14'b0000000_0000000;
		Dminus[7760] = 14'b0000000_0000000;
		Dminus[7761] = 14'b0000000_0000000;
		Dminus[7762] = 14'b0000000_0000000;
		Dminus[7763] = 14'b0000000_0000000;
		Dminus[7764] = 14'b0000000_0000000;
		Dminus[7765] = 14'b0000000_0000000;
		Dminus[7766] = 14'b0000000_0000000;
		Dminus[7767] = 14'b0000000_0000000;
		Dminus[7768] = 14'b0000000_0000000;
		Dminus[7769] = 14'b0000000_0000000;
		Dminus[7770] = 14'b0000000_0000000;
		Dminus[7771] = 14'b0000000_0000000;
		Dminus[7772] = 14'b0000000_0000000;
		Dminus[7773] = 14'b0000000_0000000;
		Dminus[7774] = 14'b0000000_0000000;
		Dminus[7775] = 14'b0000000_0000000;
		Dminus[7776] = 14'b0000000_0000000;
		Dminus[7777] = 14'b0000000_0000000;
		Dminus[7778] = 14'b0000000_0000000;
		Dminus[7779] = 14'b0000000_0000000;
		Dminus[7780] = 14'b0000000_0000000;
		Dminus[7781] = 14'b0000000_0000000;
		Dminus[7782] = 14'b0000000_0000000;
		Dminus[7783] = 14'b0000000_0000000;
		Dminus[7784] = 14'b0000000_0000000;
		Dminus[7785] = 14'b0000000_0000000;
		Dminus[7786] = 14'b0000000_0000000;
		Dminus[7787] = 14'b0000000_0000000;
		Dminus[7788] = 14'b0000000_0000000;
		Dminus[7789] = 14'b0000000_0000000;
		Dminus[7790] = 14'b0000000_0000000;
		Dminus[7791] = 14'b0000000_0000000;
		Dminus[7792] = 14'b0000000_0000000;
		Dminus[7793] = 14'b0000000_0000000;
		Dminus[7794] = 14'b0000000_0000000;
		Dminus[7795] = 14'b0000000_0000000;
		Dminus[7796] = 14'b0000000_0000000;
		Dminus[7797] = 14'b0000000_0000000;
		Dminus[7798] = 14'b0000000_0000000;
		Dminus[7799] = 14'b0000000_0000000;
		Dminus[7800] = 14'b0000000_0000000;
		Dminus[7801] = 14'b0000000_0000000;
		Dminus[7802] = 14'b0000000_0000000;
		Dminus[7803] = 14'b0000000_0000000;
		Dminus[7804] = 14'b0000000_0000000;
		Dminus[7805] = 14'b0000000_0000000;
		Dminus[7806] = 14'b0000000_0000000;
		Dminus[7807] = 14'b0000000_0000000;
		Dminus[7808] = 14'b0000000_0000000;
		Dminus[7809] = 14'b0000000_0000000;
		Dminus[7810] = 14'b0000000_0000000;
		Dminus[7811] = 14'b0000000_0000000;
		Dminus[7812] = 14'b0000000_0000000;
		Dminus[7813] = 14'b0000000_0000000;
		Dminus[7814] = 14'b0000000_0000000;
		Dminus[7815] = 14'b0000000_0000000;
		Dminus[7816] = 14'b0000000_0000000;
		Dminus[7817] = 14'b0000000_0000000;
		Dminus[7818] = 14'b0000000_0000000;
		Dminus[7819] = 14'b0000000_0000000;
		Dminus[7820] = 14'b0000000_0000000;
		Dminus[7821] = 14'b0000000_0000000;
		Dminus[7822] = 14'b0000000_0000000;
		Dminus[7823] = 14'b0000000_0000000;
		Dminus[7824] = 14'b0000000_0000000;
		Dminus[7825] = 14'b0000000_0000000;
		Dminus[7826] = 14'b0000000_0000000;
		Dminus[7827] = 14'b0000000_0000000;
		Dminus[7828] = 14'b0000000_0000000;
		Dminus[7829] = 14'b0000000_0000000;
		Dminus[7830] = 14'b0000000_0000000;
		Dminus[7831] = 14'b0000000_0000000;
		Dminus[7832] = 14'b0000000_0000000;
		Dminus[7833] = 14'b0000000_0000000;
		Dminus[7834] = 14'b0000000_0000000;
		Dminus[7835] = 14'b0000000_0000000;
		Dminus[7836] = 14'b0000000_0000000;
		Dminus[7837] = 14'b0000000_0000000;
		Dminus[7838] = 14'b0000000_0000000;
		Dminus[7839] = 14'b0000000_0000000;
		Dminus[7840] = 14'b0000000_0000000;
		Dminus[7841] = 14'b0000000_0000000;
		Dminus[7842] = 14'b0000000_0000000;
		Dminus[7843] = 14'b0000000_0000000;
		Dminus[7844] = 14'b0000000_0000000;
		Dminus[7845] = 14'b0000000_0000000;
		Dminus[7846] = 14'b0000000_0000000;
		Dminus[7847] = 14'b0000000_0000000;
		Dminus[7848] = 14'b0000000_0000000;
		Dminus[7849] = 14'b0000000_0000000;
		Dminus[7850] = 14'b0000000_0000000;
		Dminus[7851] = 14'b0000000_0000000;
		Dminus[7852] = 14'b0000000_0000000;
		Dminus[7853] = 14'b0000000_0000000;
		Dminus[7854] = 14'b0000000_0000000;
		Dminus[7855] = 14'b0000000_0000000;
		Dminus[7856] = 14'b0000000_0000000;
		Dminus[7857] = 14'b0000000_0000000;
		Dminus[7858] = 14'b0000000_0000000;
		Dminus[7859] = 14'b0000000_0000000;
		Dminus[7860] = 14'b0000000_0000000;
		Dminus[7861] = 14'b0000000_0000000;
		Dminus[7862] = 14'b0000000_0000000;
		Dminus[7863] = 14'b0000000_0000000;
		Dminus[7864] = 14'b0000000_0000000;
		Dminus[7865] = 14'b0000000_0000000;
		Dminus[7866] = 14'b0000000_0000000;
		Dminus[7867] = 14'b0000000_0000000;
		Dminus[7868] = 14'b0000000_0000000;
		Dminus[7869] = 14'b0000000_0000000;
		Dminus[7870] = 14'b0000000_0000000;
		Dminus[7871] = 14'b0000000_0000000;
		Dminus[7872] = 14'b0000000_0000000;
		Dminus[7873] = 14'b0000000_0000000;
		Dminus[7874] = 14'b0000000_0000000;
		Dminus[7875] = 14'b0000000_0000000;
		Dminus[7876] = 14'b0000000_0000000;
		Dminus[7877] = 14'b0000000_0000000;
		Dminus[7878] = 14'b0000000_0000000;
		Dminus[7879] = 14'b0000000_0000000;
		Dminus[7880] = 14'b0000000_0000000;
		Dminus[7881] = 14'b0000000_0000000;
		Dminus[7882] = 14'b0000000_0000000;
		Dminus[7883] = 14'b0000000_0000000;
		Dminus[7884] = 14'b0000000_0000000;
		Dminus[7885] = 14'b0000000_0000000;
		Dminus[7886] = 14'b0000000_0000000;
		Dminus[7887] = 14'b0000000_0000000;
		Dminus[7888] = 14'b0000000_0000000;
		Dminus[7889] = 14'b0000000_0000000;
		Dminus[7890] = 14'b0000000_0000000;
		Dminus[7891] = 14'b0000000_0000000;
		Dminus[7892] = 14'b0000000_0000000;
		Dminus[7893] = 14'b0000000_0000000;
		Dminus[7894] = 14'b0000000_0000000;
		Dminus[7895] = 14'b0000000_0000000;
		Dminus[7896] = 14'b0000000_0000000;
		Dminus[7897] = 14'b0000000_0000000;
		Dminus[7898] = 14'b0000000_0000000;
		Dminus[7899] = 14'b0000000_0000000;
		Dminus[7900] = 14'b0000000_0000000;
		Dminus[7901] = 14'b0000000_0000000;
		Dminus[7902] = 14'b0000000_0000000;
		Dminus[7903] = 14'b0000000_0000000;
		Dminus[7904] = 14'b0000000_0000000;
		Dminus[7905] = 14'b0000000_0000000;
		Dminus[7906] = 14'b0000000_0000000;
		Dminus[7907] = 14'b0000000_0000000;
		Dminus[7908] = 14'b0000000_0000000;
		Dminus[7909] = 14'b0000000_0000000;
		Dminus[7910] = 14'b0000000_0000000;
		Dminus[7911] = 14'b0000000_0000000;
		Dminus[7912] = 14'b0000000_0000000;
		Dminus[7913] = 14'b0000000_0000000;
		Dminus[7914] = 14'b0000000_0000000;
		Dminus[7915] = 14'b0000000_0000000;
		Dminus[7916] = 14'b0000000_0000000;
		Dminus[7917] = 14'b0000000_0000000;
		Dminus[7918] = 14'b0000000_0000000;
		Dminus[7919] = 14'b0000000_0000000;
		Dminus[7920] = 14'b0000000_0000000;
		Dminus[7921] = 14'b0000000_0000000;
		Dminus[7922] = 14'b0000000_0000000;
		Dminus[7923] = 14'b0000000_0000000;
		Dminus[7924] = 14'b0000000_0000000;
		Dminus[7925] = 14'b0000000_0000000;
		Dminus[7926] = 14'b0000000_0000000;
		Dminus[7927] = 14'b0000000_0000000;
		Dminus[7928] = 14'b0000000_0000000;
		Dminus[7929] = 14'b0000000_0000000;
		Dminus[7930] = 14'b0000000_0000000;
		Dminus[7931] = 14'b0000000_0000000;
		Dminus[7932] = 14'b0000000_0000000;
		Dminus[7933] = 14'b0000000_0000000;
		Dminus[7934] = 14'b0000000_0000000;
		Dminus[7935] = 14'b0000000_0000000;
		Dminus[7936] = 14'b0000000_0000000;
		Dminus[7937] = 14'b0000000_0000000;
		Dminus[7938] = 14'b0000000_0000000;
		Dminus[7939] = 14'b0000000_0000000;
		Dminus[7940] = 14'b0000000_0000000;
		Dminus[7941] = 14'b0000000_0000000;
		Dminus[7942] = 14'b0000000_0000000;
		Dminus[7943] = 14'b0000000_0000000;
		Dminus[7944] = 14'b0000000_0000000;
		Dminus[7945] = 14'b0000000_0000000;
		Dminus[7946] = 14'b0000000_0000000;
		Dminus[7947] = 14'b0000000_0000000;
		Dminus[7948] = 14'b0000000_0000000;
		Dminus[7949] = 14'b0000000_0000000;
		Dminus[7950] = 14'b0000000_0000000;
		Dminus[7951] = 14'b0000000_0000000;
		Dminus[7952] = 14'b0000000_0000000;
		Dminus[7953] = 14'b0000000_0000000;
		Dminus[7954] = 14'b0000000_0000000;
		Dminus[7955] = 14'b0000000_0000000;
		Dminus[7956] = 14'b0000000_0000000;
		Dminus[7957] = 14'b0000000_0000000;
		Dminus[7958] = 14'b0000000_0000000;
		Dminus[7959] = 14'b0000000_0000000;
		Dminus[7960] = 14'b0000000_0000000;
		Dminus[7961] = 14'b0000000_0000000;
		Dminus[7962] = 14'b0000000_0000000;
		Dminus[7963] = 14'b0000000_0000000;
		Dminus[7964] = 14'b0000000_0000000;
		Dminus[7965] = 14'b0000000_0000000;
		Dminus[7966] = 14'b0000000_0000000;
		Dminus[7967] = 14'b0000000_0000000;
		Dminus[7968] = 14'b0000000_0000000;
		Dminus[7969] = 14'b0000000_0000000;
		Dminus[7970] = 14'b0000000_0000000;
		Dminus[7971] = 14'b0000000_0000000;
		Dminus[7972] = 14'b0000000_0000000;
		Dminus[7973] = 14'b0000000_0000000;
		Dminus[7974] = 14'b0000000_0000000;
		Dminus[7975] = 14'b0000000_0000000;
		Dminus[7976] = 14'b0000000_0000000;
		Dminus[7977] = 14'b0000000_0000000;
		Dminus[7978] = 14'b0000000_0000000;
		Dminus[7979] = 14'b0000000_0000000;
		Dminus[7980] = 14'b0000000_0000000;
		Dminus[7981] = 14'b0000000_0000000;
		Dminus[7982] = 14'b0000000_0000000;
		Dminus[7983] = 14'b0000000_0000000;
		Dminus[7984] = 14'b0000000_0000000;
		Dminus[7985] = 14'b0000000_0000000;
		Dminus[7986] = 14'b0000000_0000000;
		Dminus[7987] = 14'b0000000_0000000;
		Dminus[7988] = 14'b0000000_0000000;
		Dminus[7989] = 14'b0000000_0000000;
		Dminus[7990] = 14'b0000000_0000000;
		Dminus[7991] = 14'b0000000_0000000;
		Dminus[7992] = 14'b0000000_0000000;
		Dminus[7993] = 14'b0000000_0000000;
		Dminus[7994] = 14'b0000000_0000000;
		Dminus[7995] = 14'b0000000_0000000;
		Dminus[7996] = 14'b0000000_0000000;
		Dminus[7997] = 14'b0000000_0000000;
		Dminus[7998] = 14'b0000000_0000000;
		Dminus[7999] = 14'b0000000_0000000;
		Dminus[8000] = 14'b0000000_0000000;
		Dminus[8001] = 14'b0000000_0000000;
		Dminus[8002] = 14'b0000000_0000000;
		Dminus[8003] = 14'b0000000_0000000;
		Dminus[8004] = 14'b0000000_0000000;
		Dminus[8005] = 14'b0000000_0000000;
		Dminus[8006] = 14'b0000000_0000000;
		Dminus[8007] = 14'b0000000_0000000;
		Dminus[8008] = 14'b0000000_0000000;
		Dminus[8009] = 14'b0000000_0000000;
		Dminus[8010] = 14'b0000000_0000000;
		Dminus[8011] = 14'b0000000_0000000;
		Dminus[8012] = 14'b0000000_0000000;
		Dminus[8013] = 14'b0000000_0000000;
		Dminus[8014] = 14'b0000000_0000000;
		Dminus[8015] = 14'b0000000_0000000;
		Dminus[8016] = 14'b0000000_0000000;
		Dminus[8017] = 14'b0000000_0000000;
		Dminus[8018] = 14'b0000000_0000000;
		Dminus[8019] = 14'b0000000_0000000;
		Dminus[8020] = 14'b0000000_0000000;
		Dminus[8021] = 14'b0000000_0000000;
		Dminus[8022] = 14'b0000000_0000000;
		Dminus[8023] = 14'b0000000_0000000;
		Dminus[8024] = 14'b0000000_0000000;
		Dminus[8025] = 14'b0000000_0000000;
		Dminus[8026] = 14'b0000000_0000000;
		Dminus[8027] = 14'b0000000_0000000;
		Dminus[8028] = 14'b0000000_0000000;
		Dminus[8029] = 14'b0000000_0000000;
		Dminus[8030] = 14'b0000000_0000000;
		Dminus[8031] = 14'b0000000_0000000;
		Dminus[8032] = 14'b0000000_0000000;
		Dminus[8033] = 14'b0000000_0000000;
		Dminus[8034] = 14'b0000000_0000000;
		Dminus[8035] = 14'b0000000_0000000;
		Dminus[8036] = 14'b0000000_0000000;
		Dminus[8037] = 14'b0000000_0000000;
		Dminus[8038] = 14'b0000000_0000000;
		Dminus[8039] = 14'b0000000_0000000;
		Dminus[8040] = 14'b0000000_0000000;
		Dminus[8041] = 14'b0000000_0000000;
		Dminus[8042] = 14'b0000000_0000000;
		Dminus[8043] = 14'b0000000_0000000;
		Dminus[8044] = 14'b0000000_0000000;
		Dminus[8045] = 14'b0000000_0000000;
		Dminus[8046] = 14'b0000000_0000000;
		Dminus[8047] = 14'b0000000_0000000;
		Dminus[8048] = 14'b0000000_0000000;
		Dminus[8049] = 14'b0000000_0000000;
		Dminus[8050] = 14'b0000000_0000000;
		Dminus[8051] = 14'b0000000_0000000;
		Dminus[8052] = 14'b0000000_0000000;
		Dminus[8053] = 14'b0000000_0000000;
		Dminus[8054] = 14'b0000000_0000000;
		Dminus[8055] = 14'b0000000_0000000;
		Dminus[8056] = 14'b0000000_0000000;
		Dminus[8057] = 14'b0000000_0000000;
		Dminus[8058] = 14'b0000000_0000000;
		Dminus[8059] = 14'b0000000_0000000;
		Dminus[8060] = 14'b0000000_0000000;
		Dminus[8061] = 14'b0000000_0000000;
		Dminus[8062] = 14'b0000000_0000000;
		Dminus[8063] = 14'b0000000_0000000;
		Dminus[8064] = 14'b0000000_0000000;
		Dminus[8065] = 14'b0000000_0000000;
		Dminus[8066] = 14'b0000000_0000000;
		Dminus[8067] = 14'b0000000_0000000;
		Dminus[8068] = 14'b0000000_0000000;
		Dminus[8069] = 14'b0000000_0000000;
		Dminus[8070] = 14'b0000000_0000000;
		Dminus[8071] = 14'b0000000_0000000;
		Dminus[8072] = 14'b0000000_0000000;
		Dminus[8073] = 14'b0000000_0000000;
		Dminus[8074] = 14'b0000000_0000000;
		Dminus[8075] = 14'b0000000_0000000;
		Dminus[8076] = 14'b0000000_0000000;
		Dminus[8077] = 14'b0000000_0000000;
		Dminus[8078] = 14'b0000000_0000000;
		Dminus[8079] = 14'b0000000_0000000;
		Dminus[8080] = 14'b0000000_0000000;
		Dminus[8081] = 14'b0000000_0000000;
		Dminus[8082] = 14'b0000000_0000000;
		Dminus[8083] = 14'b0000000_0000000;
		Dminus[8084] = 14'b0000000_0000000;
		Dminus[8085] = 14'b0000000_0000000;
		Dminus[8086] = 14'b0000000_0000000;
		Dminus[8087] = 14'b0000000_0000000;
		Dminus[8088] = 14'b0000000_0000000;
		Dminus[8089] = 14'b0000000_0000000;
		Dminus[8090] = 14'b0000000_0000000;
		Dminus[8091] = 14'b0000000_0000000;
		Dminus[8092] = 14'b0000000_0000000;
		Dminus[8093] = 14'b0000000_0000000;
		Dminus[8094] = 14'b0000000_0000000;
		Dminus[8095] = 14'b0000000_0000000;
		Dminus[8096] = 14'b0000000_0000000;
		Dminus[8097] = 14'b0000000_0000000;
		Dminus[8098] = 14'b0000000_0000000;
		Dminus[8099] = 14'b0000000_0000000;
		Dminus[8100] = 14'b0000000_0000000;
		Dminus[8101] = 14'b0000000_0000000;
		Dminus[8102] = 14'b0000000_0000000;
		Dminus[8103] = 14'b0000000_0000000;
		Dminus[8104] = 14'b0000000_0000000;
		Dminus[8105] = 14'b0000000_0000000;
		Dminus[8106] = 14'b0000000_0000000;
		Dminus[8107] = 14'b0000000_0000000;
		Dminus[8108] = 14'b0000000_0000000;
		Dminus[8109] = 14'b0000000_0000000;
		Dminus[8110] = 14'b0000000_0000000;
		Dminus[8111] = 14'b0000000_0000000;
		Dminus[8112] = 14'b0000000_0000000;
		Dminus[8113] = 14'b0000000_0000000;
		Dminus[8114] = 14'b0000000_0000000;
		Dminus[8115] = 14'b0000000_0000000;
		Dminus[8116] = 14'b0000000_0000000;
		Dminus[8117] = 14'b0000000_0000000;
		Dminus[8118] = 14'b0000000_0000000;
		Dminus[8119] = 14'b0000000_0000000;
		Dminus[8120] = 14'b0000000_0000000;
		Dminus[8121] = 14'b0000000_0000000;
		Dminus[8122] = 14'b0000000_0000000;
		Dminus[8123] = 14'b0000000_0000000;
		Dminus[8124] = 14'b0000000_0000000;
		Dminus[8125] = 14'b0000000_0000000;
		Dminus[8126] = 14'b0000000_0000000;
		Dminus[8127] = 14'b0000000_0000000;
		Dminus[8128] = 14'b0000000_0000000;
		Dminus[8129] = 14'b0000000_0000000;
		Dminus[8130] = 14'b0000000_0000000;
		Dminus[8131] = 14'b0000000_0000000;
		Dminus[8132] = 14'b0000000_0000000;
		Dminus[8133] = 14'b0000000_0000000;
		Dminus[8134] = 14'b0000000_0000000;
		Dminus[8135] = 14'b0000000_0000000;
		Dminus[8136] = 14'b0000000_0000000;
		Dminus[8137] = 14'b0000000_0000000;
		Dminus[8138] = 14'b0000000_0000000;
		Dminus[8139] = 14'b0000000_0000000;
		Dminus[8140] = 14'b0000000_0000000;
		Dminus[8141] = 14'b0000000_0000000;
		Dminus[8142] = 14'b0000000_0000000;
		Dminus[8143] = 14'b0000000_0000000;
		Dminus[8144] = 14'b0000000_0000000;
		Dminus[8145] = 14'b0000000_0000000;
		Dminus[8146] = 14'b0000000_0000000;
		Dminus[8147] = 14'b0000000_0000000;
		Dminus[8148] = 14'b0000000_0000000;
		Dminus[8149] = 14'b0000000_0000000;
		Dminus[8150] = 14'b0000000_0000000;
		Dminus[8151] = 14'b0000000_0000000;
		Dminus[8152] = 14'b0000000_0000000;
		Dminus[8153] = 14'b0000000_0000000;
		Dminus[8154] = 14'b0000000_0000000;
		Dminus[8155] = 14'b0000000_0000000;
		Dminus[8156] = 14'b0000000_0000000;
		Dminus[8157] = 14'b0000000_0000000;
		Dminus[8158] = 14'b0000000_0000000;
		Dminus[8159] = 14'b0000000_0000000;
		Dminus[8160] = 14'b0000000_0000000;
		Dminus[8161] = 14'b0000000_0000000;
		Dminus[8162] = 14'b0000000_0000000;
		Dminus[8163] = 14'b0000000_0000000;
		Dminus[8164] = 14'b0000000_0000000;
		Dminus[8165] = 14'b0000000_0000000;
		Dminus[8166] = 14'b0000000_0000000;
		Dminus[8167] = 14'b0000000_0000000;
		Dminus[8168] = 14'b0000000_0000000;
		Dminus[8169] = 14'b0000000_0000000;
		Dminus[8170] = 14'b0000000_0000000;
		Dminus[8171] = 14'b0000000_0000000;
		Dminus[8172] = 14'b0000000_0000000;
		Dminus[8173] = 14'b0000000_0000000;
		Dminus[8174] = 14'b0000000_0000000;
		Dminus[8175] = 14'b0000000_0000000;
		Dminus[8176] = 14'b0000000_0000000;
		Dminus[8177] = 14'b0000000_0000000;
		Dminus[8178] = 14'b0000000_0000000;
		Dminus[8179] = 14'b0000000_0000000;
		Dminus[8180] = 14'b0000000_0000000;
		Dminus[8181] = 14'b0000000_0000000;
		Dminus[8182] = 14'b0000000_0000000;
		Dminus[8183] = 14'b0000000_0000000;
		Dminus[8184] = 14'b0000000_0000000;
		Dminus[8185] = 14'b0000000_0000000;
		Dminus[8186] = 14'b0000000_0000000;
		Dminus[8187] = 14'b0000000_0000000;
		Dminus[8188] = 14'b0000000_0000000;
		Dminus[8189] = 14'b0000000_0000000;
		Dminus[8190] = 14'b0000000_0000000;
		Dminus[8191] = 14'b0000000_0000000;
		Dplus[1] = 14'b0000001_0000000;
		Dplus[2] = 14'b0000000_1111111;
		Dplus[3] = 14'b0000000_1111111;
		Dplus[4] = 14'b0000000_1111110;
		Dplus[5] = 14'b0000000_1111110;
		Dplus[6] = 14'b0000000_1111101;
		Dplus[7] = 14'b0000000_1111101;
		Dplus[8] = 14'b0000000_1111100;
		Dplus[9] = 14'b0000000_1111100;
		Dplus[10] = 14'b0000000_1111011;
		Dplus[11] = 14'b0000000_1111011;
		Dplus[12] = 14'b0000000_1111010;
		Dplus[13] = 14'b0000000_1111010;
		Dplus[14] = 14'b0000000_1111001;
		Dplus[15] = 14'b0000000_1111001;
		Dplus[16] = 14'b0000000_1111000;
		Dplus[17] = 14'b0000000_1111000;
		Dplus[18] = 14'b0000000_1110111;
		Dplus[19] = 14'b0000000_1110111;
		Dplus[20] = 14'b0000000_1110110;
		Dplus[21] = 14'b0000000_1110110;
		Dplus[22] = 14'b0000000_1110101;
		Dplus[23] = 14'b0000000_1110101;
		Dplus[24] = 14'b0000000_1110100;
		Dplus[25] = 14'b0000000_1110100;
		Dplus[26] = 14'b0000000_1110011;
		Dplus[27] = 14'b0000000_1110011;
		Dplus[28] = 14'b0000000_1110011;
		Dplus[29] = 14'b0000000_1110010;
		Dplus[30] = 14'b0000000_1110010;
		Dplus[31] = 14'b0000000_1110001;
		Dplus[32] = 14'b0000000_1110001;
		Dplus[33] = 14'b0000000_1110000;
		Dplus[34] = 14'b0000000_1110000;
		Dplus[35] = 14'b0000000_1101111;
		Dplus[36] = 14'b0000000_1101111;
		Dplus[37] = 14'b0000000_1101110;
		Dplus[38] = 14'b0000000_1101110;
		Dplus[39] = 14'b0000000_1101110;
		Dplus[40] = 14'b0000000_1101101;
		Dplus[41] = 14'b0000000_1101101;
		Dplus[42] = 14'b0000000_1101100;
		Dplus[43] = 14'b0000000_1101100;
		Dplus[44] = 14'b0000000_1101011;
		Dplus[45] = 14'b0000000_1101011;
		Dplus[46] = 14'b0000000_1101010;
		Dplus[47] = 14'b0000000_1101010;
		Dplus[48] = 14'b0000000_1101010;
		Dplus[49] = 14'b0000000_1101001;
		Dplus[50] = 14'b0000000_1101001;
		Dplus[51] = 14'b0000000_1101000;
		Dplus[52] = 14'b0000000_1101000;
		Dplus[53] = 14'b0000000_1100111;
		Dplus[54] = 14'b0000000_1100111;
		Dplus[55] = 14'b0000000_1100111;
		Dplus[56] = 14'b0000000_1100110;
		Dplus[57] = 14'b0000000_1100110;
		Dplus[58] = 14'b0000000_1100101;
		Dplus[59] = 14'b0000000_1100101;
		Dplus[60] = 14'b0000000_1100100;
		Dplus[61] = 14'b0000000_1100100;
		Dplus[62] = 14'b0000000_1100100;
		Dplus[63] = 14'b0000000_1100011;
		Dplus[64] = 14'b0000000_1100011;
		Dplus[65] = 14'b0000000_1100010;
		Dplus[66] = 14'b0000000_1100010;
		Dplus[67] = 14'b0000000_1100010;
		Dplus[68] = 14'b0000000_1100001;
		Dplus[69] = 14'b0000000_1100001;
		Dplus[70] = 14'b0000000_1100000;
		Dplus[71] = 14'b0000000_1100000;
		Dplus[72] = 14'b0000000_1011111;
		Dplus[73] = 14'b0000000_1011111;
		Dplus[74] = 14'b0000000_1011111;
		Dplus[75] = 14'b0000000_1011110;
		Dplus[76] = 14'b0000000_1011110;
		Dplus[77] = 14'b0000000_1011101;
		Dplus[78] = 14'b0000000_1011101;
		Dplus[79] = 14'b0000000_1011101;
		Dplus[80] = 14'b0000000_1011100;
		Dplus[81] = 14'b0000000_1011100;
		Dplus[82] = 14'b0000000_1011100;
		Dplus[83] = 14'b0000000_1011011;
		Dplus[84] = 14'b0000000_1011011;
		Dplus[85] = 14'b0000000_1011010;
		Dplus[86] = 14'b0000000_1011010;
		Dplus[87] = 14'b0000000_1011010;
		Dplus[88] = 14'b0000000_1011001;
		Dplus[89] = 14'b0000000_1011001;
		Dplus[90] = 14'b0000000_1011000;
		Dplus[91] = 14'b0000000_1011000;
		Dplus[92] = 14'b0000000_1011000;
		Dplus[93] = 14'b0000000_1010111;
		Dplus[94] = 14'b0000000_1010111;
		Dplus[95] = 14'b0000000_1010111;
		Dplus[96] = 14'b0000000_1010110;
		Dplus[97] = 14'b0000000_1010110;
		Dplus[98] = 14'b0000000_1010101;
		Dplus[99] = 14'b0000000_1010101;
		Dplus[100] = 14'b0000000_1010101;
		Dplus[101] = 14'b0000000_1010100;
		Dplus[102] = 14'b0000000_1010100;
		Dplus[103] = 14'b0000000_1010100;
		Dplus[104] = 14'b0000000_1010011;
		Dplus[105] = 14'b0000000_1010011;
		Dplus[106] = 14'b0000000_1010011;
		Dplus[107] = 14'b0000000_1010010;
		Dplus[108] = 14'b0000000_1010010;
		Dplus[109] = 14'b0000000_1010001;
		Dplus[110] = 14'b0000000_1010001;
		Dplus[111] = 14'b0000000_1010001;
		Dplus[112] = 14'b0000000_1010000;
		Dplus[113] = 14'b0000000_1010000;
		Dplus[114] = 14'b0000000_1010000;
		Dplus[115] = 14'b0000000_1001111;
		Dplus[116] = 14'b0000000_1001111;
		Dplus[117] = 14'b0000000_1001111;
		Dplus[118] = 14'b0000000_1001110;
		Dplus[119] = 14'b0000000_1001110;
		Dplus[120] = 14'b0000000_1001110;
		Dplus[121] = 14'b0000000_1001101;
		Dplus[122] = 14'b0000000_1001101;
		Dplus[123] = 14'b0000000_1001101;
		Dplus[124] = 14'b0000000_1001100;
		Dplus[125] = 14'b0000000_1001100;
		Dplus[126] = 14'b0000000_1001100;
		Dplus[127] = 14'b0000000_1001011;
		Dplus[128] = 14'b0000000_1001011;
		Dplus[129] = 14'b0000000_1001011;
		Dplus[130] = 14'b0000000_1001010;
		Dplus[131] = 14'b0000000_1001010;
		Dplus[132] = 14'b0000000_1001010;
		Dplus[133] = 14'b0000000_1001001;
		Dplus[134] = 14'b0000000_1001001;
		Dplus[135] = 14'b0000000_1001001;
		Dplus[136] = 14'b0000000_1001000;
		Dplus[137] = 14'b0000000_1001000;
		Dplus[138] = 14'b0000000_1001000;
		Dplus[139] = 14'b0000000_1000111;
		Dplus[140] = 14'b0000000_1000111;
		Dplus[141] = 14'b0000000_1000111;
		Dplus[142] = 14'b0000000_1000110;
		Dplus[143] = 14'b0000000_1000110;
		Dplus[144] = 14'b0000000_1000110;
		Dplus[145] = 14'b0000000_1000101;
		Dplus[146] = 14'b0000000_1000101;
		Dplus[147] = 14'b0000000_1000101;
		Dplus[148] = 14'b0000000_1000100;
		Dplus[149] = 14'b0000000_1000100;
		Dplus[150] = 14'b0000000_1000100;
		Dplus[151] = 14'b0000000_1000100;
		Dplus[152] = 14'b0000000_1000011;
		Dplus[153] = 14'b0000000_1000011;
		Dplus[154] = 14'b0000000_1000011;
		Dplus[155] = 14'b0000000_1000010;
		Dplus[156] = 14'b0000000_1000010;
		Dplus[157] = 14'b0000000_1000010;
		Dplus[158] = 14'b0000000_1000001;
		Dplus[159] = 14'b0000000_1000001;
		Dplus[160] = 14'b0000000_1000001;
		Dplus[161] = 14'b0000000_1000001;
		Dplus[162] = 14'b0000000_1000000;
		Dplus[163] = 14'b0000000_1000000;
		Dplus[164] = 14'b0000000_1000000;
		Dplus[165] = 14'b0000000_0111111;
		Dplus[166] = 14'b0000000_0111111;
		Dplus[167] = 14'b0000000_0111111;
		Dplus[168] = 14'b0000000_0111110;
		Dplus[169] = 14'b0000000_0111110;
		Dplus[170] = 14'b0000000_0111110;
		Dplus[171] = 14'b0000000_0111110;
		Dplus[172] = 14'b0000000_0111101;
		Dplus[173] = 14'b0000000_0111101;
		Dplus[174] = 14'b0000000_0111101;
		Dplus[175] = 14'b0000000_0111100;
		Dplus[176] = 14'b0000000_0111100;
		Dplus[177] = 14'b0000000_0111100;
		Dplus[178] = 14'b0000000_0111100;
		Dplus[179] = 14'b0000000_0111011;
		Dplus[180] = 14'b0000000_0111011;
		Dplus[181] = 14'b0000000_0111011;
		Dplus[182] = 14'b0000000_0111011;
		Dplus[183] = 14'b0000000_0111010;
		Dplus[184] = 14'b0000000_0111010;
		Dplus[185] = 14'b0000000_0111010;
		Dplus[186] = 14'b0000000_0111001;
		Dplus[187] = 14'b0000000_0111001;
		Dplus[188] = 14'b0000000_0111001;
		Dplus[189] = 14'b0000000_0111001;
		Dplus[190] = 14'b0000000_0111000;
		Dplus[191] = 14'b0000000_0111000;
		Dplus[192] = 14'b0000000_0111000;
		Dplus[193] = 14'b0000000_0111000;
		Dplus[194] = 14'b0000000_0110111;
		Dplus[195] = 14'b0000000_0110111;
		Dplus[196] = 14'b0000000_0110111;
		Dplus[197] = 14'b0000000_0110111;
		Dplus[198] = 14'b0000000_0110110;
		Dplus[199] = 14'b0000000_0110110;
		Dplus[200] = 14'b0000000_0110110;
		Dplus[201] = 14'b0000000_0110110;
		Dplus[202] = 14'b0000000_0110101;
		Dplus[203] = 14'b0000000_0110101;
		Dplus[204] = 14'b0000000_0110101;
		Dplus[205] = 14'b0000000_0110101;
		Dplus[206] = 14'b0000000_0110100;
		Dplus[207] = 14'b0000000_0110100;
		Dplus[208] = 14'b0000000_0110100;
		Dplus[209] = 14'b0000000_0110100;
		Dplus[210] = 14'b0000000_0110011;
		Dplus[211] = 14'b0000000_0110011;
		Dplus[212] = 14'b0000000_0110011;
		Dplus[213] = 14'b0000000_0110011;
		Dplus[214] = 14'b0000000_0110010;
		Dplus[215] = 14'b0000000_0110010;
		Dplus[216] = 14'b0000000_0110010;
		Dplus[217] = 14'b0000000_0110010;
		Dplus[218] = 14'b0000000_0110001;
		Dplus[219] = 14'b0000000_0110001;
		Dplus[220] = 14'b0000000_0110001;
		Dplus[221] = 14'b0000000_0110001;
		Dplus[222] = 14'b0000000_0110001;
		Dplus[223] = 14'b0000000_0110000;
		Dplus[224] = 14'b0000000_0110000;
		Dplus[225] = 14'b0000000_0110000;
		Dplus[226] = 14'b0000000_0110000;
		Dplus[227] = 14'b0000000_0101111;
		Dplus[228] = 14'b0000000_0101111;
		Dplus[229] = 14'b0000000_0101111;
		Dplus[230] = 14'b0000000_0101111;
		Dplus[231] = 14'b0000000_0101110;
		Dplus[232] = 14'b0000000_0101110;
		Dplus[233] = 14'b0000000_0101110;
		Dplus[234] = 14'b0000000_0101110;
		Dplus[235] = 14'b0000000_0101110;
		Dplus[236] = 14'b0000000_0101101;
		Dplus[237] = 14'b0000000_0101101;
		Dplus[238] = 14'b0000000_0101101;
		Dplus[239] = 14'b0000000_0101101;
		Dplus[240] = 14'b0000000_0101101;
		Dplus[241] = 14'b0000000_0101100;
		Dplus[242] = 14'b0000000_0101100;
		Dplus[243] = 14'b0000000_0101100;
		Dplus[244] = 14'b0000000_0101100;
		Dplus[245] = 14'b0000000_0101011;
		Dplus[246] = 14'b0000000_0101011;
		Dplus[247] = 14'b0000000_0101011;
		Dplus[248] = 14'b0000000_0101011;
		Dplus[249] = 14'b0000000_0101011;
		Dplus[250] = 14'b0000000_0101010;
		Dplus[251] = 14'b0000000_0101010;
		Dplus[252] = 14'b0000000_0101010;
		Dplus[253] = 14'b0000000_0101010;
		Dplus[254] = 14'b0000000_0101010;
		Dplus[255] = 14'b0000000_0101001;
		Dplus[256] = 14'b0000000_0101001;
		Dplus[257] = 14'b0000000_0101001;
		Dplus[258] = 14'b0000000_0101001;
		Dplus[259] = 14'b0000000_0101001;
		Dplus[260] = 14'b0000000_0101000;
		Dplus[261] = 14'b0000000_0101000;
		Dplus[262] = 14'b0000000_0101000;
		Dplus[263] = 14'b0000000_0101000;
		Dplus[264] = 14'b0000000_0101000;
		Dplus[265] = 14'b0000000_0100111;
		Dplus[266] = 14'b0000000_0100111;
		Dplus[267] = 14'b0000000_0100111;
		Dplus[268] = 14'b0000000_0100111;
		Dplus[269] = 14'b0000000_0100111;
		Dplus[270] = 14'b0000000_0100110;
		Dplus[271] = 14'b0000000_0100110;
		Dplus[272] = 14'b0000000_0100110;
		Dplus[273] = 14'b0000000_0100110;
		Dplus[274] = 14'b0000000_0100110;
		Dplus[275] = 14'b0000000_0100110;
		Dplus[276] = 14'b0000000_0100101;
		Dplus[277] = 14'b0000000_0100101;
		Dplus[278] = 14'b0000000_0100101;
		Dplus[279] = 14'b0000000_0100101;
		Dplus[280] = 14'b0000000_0100101;
		Dplus[281] = 14'b0000000_0100100;
		Dplus[282] = 14'b0000000_0100100;
		Dplus[283] = 14'b0000000_0100100;
		Dplus[284] = 14'b0000000_0100100;
		Dplus[285] = 14'b0000000_0100100;
		Dplus[286] = 14'b0000000_0100100;
		Dplus[287] = 14'b0000000_0100011;
		Dplus[288] = 14'b0000000_0100011;
		Dplus[289] = 14'b0000000_0100011;
		Dplus[290] = 14'b0000000_0100011;
		Dplus[291] = 14'b0000000_0100011;
		Dplus[292] = 14'b0000000_0100011;
		Dplus[293] = 14'b0000000_0100010;
		Dplus[294] = 14'b0000000_0100010;
		Dplus[295] = 14'b0000000_0100010;
		Dplus[296] = 14'b0000000_0100010;
		Dplus[297] = 14'b0000000_0100010;
		Dplus[298] = 14'b0000000_0100010;
		Dplus[299] = 14'b0000000_0100001;
		Dplus[300] = 14'b0000000_0100001;
		Dplus[301] = 14'b0000000_0100001;
		Dplus[302] = 14'b0000000_0100001;
		Dplus[303] = 14'b0000000_0100001;
		Dplus[304] = 14'b0000000_0100001;
		Dplus[305] = 14'b0000000_0100000;
		Dplus[306] = 14'b0000000_0100000;
		Dplus[307] = 14'b0000000_0100000;
		Dplus[308] = 14'b0000000_0100000;
		Dplus[309] = 14'b0000000_0100000;
		Dplus[310] = 14'b0000000_0100000;
		Dplus[311] = 14'b0000000_0011111;
		Dplus[312] = 14'b0000000_0011111;
		Dplus[313] = 14'b0000000_0011111;
		Dplus[314] = 14'b0000000_0011111;
		Dplus[315] = 14'b0000000_0011111;
		Dplus[316] = 14'b0000000_0011111;
		Dplus[317] = 14'b0000000_0011111;
		Dplus[318] = 14'b0000000_0011110;
		Dplus[319] = 14'b0000000_0011110;
		Dplus[320] = 14'b0000000_0011110;
		Dplus[321] = 14'b0000000_0011110;
		Dplus[322] = 14'b0000000_0011110;
		Dplus[323] = 14'b0000000_0011110;
		Dplus[324] = 14'b0000000_0011101;
		Dplus[325] = 14'b0000000_0011101;
		Dplus[326] = 14'b0000000_0011101;
		Dplus[327] = 14'b0000000_0011101;
		Dplus[328] = 14'b0000000_0011101;
		Dplus[329] = 14'b0000000_0011101;
		Dplus[330] = 14'b0000000_0011101;
		Dplus[331] = 14'b0000000_0011100;
		Dplus[332] = 14'b0000000_0011100;
		Dplus[333] = 14'b0000000_0011100;
		Dplus[334] = 14'b0000000_0011100;
		Dplus[335] = 14'b0000000_0011100;
		Dplus[336] = 14'b0000000_0011100;
		Dplus[337] = 14'b0000000_0011100;
		Dplus[338] = 14'b0000000_0011011;
		Dplus[339] = 14'b0000000_0011011;
		Dplus[340] = 14'b0000000_0011011;
		Dplus[341] = 14'b0000000_0011011;
		Dplus[342] = 14'b0000000_0011011;
		Dplus[343] = 14'b0000000_0011011;
		Dplus[344] = 14'b0000000_0011011;
		Dplus[345] = 14'b0000000_0011011;
		Dplus[346] = 14'b0000000_0011010;
		Dplus[347] = 14'b0000000_0011010;
		Dplus[348] = 14'b0000000_0011010;
		Dplus[349] = 14'b0000000_0011010;
		Dplus[350] = 14'b0000000_0011010;
		Dplus[351] = 14'b0000000_0011010;
		Dplus[352] = 14'b0000000_0011010;
		Dplus[353] = 14'b0000000_0011001;
		Dplus[354] = 14'b0000000_0011001;
		Dplus[355] = 14'b0000000_0011001;
		Dplus[356] = 14'b0000000_0011001;
		Dplus[357] = 14'b0000000_0011001;
		Dplus[358] = 14'b0000000_0011001;
		Dplus[359] = 14'b0000000_0011001;
		Dplus[360] = 14'b0000000_0011001;
		Dplus[361] = 14'b0000000_0011000;
		Dplus[362] = 14'b0000000_0011000;
		Dplus[363] = 14'b0000000_0011000;
		Dplus[364] = 14'b0000000_0011000;
		Dplus[365] = 14'b0000000_0011000;
		Dplus[366] = 14'b0000000_0011000;
		Dplus[367] = 14'b0000000_0011000;
		Dplus[368] = 14'b0000000_0011000;
		Dplus[369] = 14'b0000000_0010111;
		Dplus[370] = 14'b0000000_0010111;
		Dplus[371] = 14'b0000000_0010111;
		Dplus[372] = 14'b0000000_0010111;
		Dplus[373] = 14'b0000000_0010111;
		Dplus[374] = 14'b0000000_0010111;
		Dplus[375] = 14'b0000000_0010111;
		Dplus[376] = 14'b0000000_0010111;
		Dplus[377] = 14'b0000000_0010111;
		Dplus[378] = 14'b0000000_0010110;
		Dplus[379] = 14'b0000000_0010110;
		Dplus[380] = 14'b0000000_0010110;
		Dplus[381] = 14'b0000000_0010110;
		Dplus[382] = 14'b0000000_0010110;
		Dplus[383] = 14'b0000000_0010110;
		Dplus[384] = 14'b0000000_0010110;
		Dplus[385] = 14'b0000000_0010110;
		Dplus[386] = 14'b0000000_0010110;
		Dplus[387] = 14'b0000000_0010101;
		Dplus[388] = 14'b0000000_0010101;
		Dplus[389] = 14'b0000000_0010101;
		Dplus[390] = 14'b0000000_0010101;
		Dplus[391] = 14'b0000000_0010101;
		Dplus[392] = 14'b0000000_0010101;
		Dplus[393] = 14'b0000000_0010101;
		Dplus[394] = 14'b0000000_0010101;
		Dplus[395] = 14'b0000000_0010101;
		Dplus[396] = 14'b0000000_0010100;
		Dplus[397] = 14'b0000000_0010100;
		Dplus[398] = 14'b0000000_0010100;
		Dplus[399] = 14'b0000000_0010100;
		Dplus[400] = 14'b0000000_0010100;
		Dplus[401] = 14'b0000000_0010100;
		Dplus[402] = 14'b0000000_0010100;
		Dplus[403] = 14'b0000000_0010100;
		Dplus[404] = 14'b0000000_0010100;
		Dplus[405] = 14'b0000000_0010100;
		Dplus[406] = 14'b0000000_0010011;
		Dplus[407] = 14'b0000000_0010011;
		Dplus[408] = 14'b0000000_0010011;
		Dplus[409] = 14'b0000000_0010011;
		Dplus[410] = 14'b0000000_0010011;
		Dplus[411] = 14'b0000000_0010011;
		Dplus[412] = 14'b0000000_0010011;
		Dplus[413] = 14'b0000000_0010011;
		Dplus[414] = 14'b0000000_0010011;
		Dplus[415] = 14'b0000000_0010011;
		Dplus[416] = 14'b0000000_0010010;
		Dplus[417] = 14'b0000000_0010010;
		Dplus[418] = 14'b0000000_0010010;
		Dplus[419] = 14'b0000000_0010010;
		Dplus[420] = 14'b0000000_0010010;
		Dplus[421] = 14'b0000000_0010010;
		Dplus[422] = 14'b0000000_0010010;
		Dplus[423] = 14'b0000000_0010010;
		Dplus[424] = 14'b0000000_0010010;
		Dplus[425] = 14'b0000000_0010010;
		Dplus[426] = 14'b0000000_0010010;
		Dplus[427] = 14'b0000000_0010001;
		Dplus[428] = 14'b0000000_0010001;
		Dplus[429] = 14'b0000000_0010001;
		Dplus[430] = 14'b0000000_0010001;
		Dplus[431] = 14'b0000000_0010001;
		Dplus[432] = 14'b0000000_0010001;
		Dplus[433] = 14'b0000000_0010001;
		Dplus[434] = 14'b0000000_0010001;
		Dplus[435] = 14'b0000000_0010001;
		Dplus[436] = 14'b0000000_0010001;
		Dplus[437] = 14'b0000000_0010001;
		Dplus[438] = 14'b0000000_0010000;
		Dplus[439] = 14'b0000000_0010000;
		Dplus[440] = 14'b0000000_0010000;
		Dplus[441] = 14'b0000000_0010000;
		Dplus[442] = 14'b0000000_0010000;
		Dplus[443] = 14'b0000000_0010000;
		Dplus[444] = 14'b0000000_0010000;
		Dplus[445] = 14'b0000000_0010000;
		Dplus[446] = 14'b0000000_0010000;
		Dplus[447] = 14'b0000000_0010000;
		Dplus[448] = 14'b0000000_0010000;
		Dplus[449] = 14'b0000000_0010000;
		Dplus[450] = 14'b0000000_0001111;
		Dplus[451] = 14'b0000000_0001111;
		Dplus[452] = 14'b0000000_0001111;
		Dplus[453] = 14'b0000000_0001111;
		Dplus[454] = 14'b0000000_0001111;
		Dplus[455] = 14'b0000000_0001111;
		Dplus[456] = 14'b0000000_0001111;
		Dplus[457] = 14'b0000000_0001111;
		Dplus[458] = 14'b0000000_0001111;
		Dplus[459] = 14'b0000000_0001111;
		Dplus[460] = 14'b0000000_0001111;
		Dplus[461] = 14'b0000000_0001111;
		Dplus[462] = 14'b0000000_0001111;
		Dplus[463] = 14'b0000000_0001110;
		Dplus[464] = 14'b0000000_0001110;
		Dplus[465] = 14'b0000000_0001110;
		Dplus[466] = 14'b0000000_0001110;
		Dplus[467] = 14'b0000000_0001110;
		Dplus[468] = 14'b0000000_0001110;
		Dplus[469] = 14'b0000000_0001110;
		Dplus[470] = 14'b0000000_0001110;
		Dplus[471] = 14'b0000000_0001110;
		Dplus[472] = 14'b0000000_0001110;
		Dplus[473] = 14'b0000000_0001110;
		Dplus[474] = 14'b0000000_0001110;
		Dplus[475] = 14'b0000000_0001110;
		Dplus[476] = 14'b0000000_0001110;
		Dplus[477] = 14'b0000000_0001101;
		Dplus[478] = 14'b0000000_0001101;
		Dplus[479] = 14'b0000000_0001101;
		Dplus[480] = 14'b0000000_0001101;
		Dplus[481] = 14'b0000000_0001101;
		Dplus[482] = 14'b0000000_0001101;
		Dplus[483] = 14'b0000000_0001101;
		Dplus[484] = 14'b0000000_0001101;
		Dplus[485] = 14'b0000000_0001101;
		Dplus[486] = 14'b0000000_0001101;
		Dplus[487] = 14'b0000000_0001101;
		Dplus[488] = 14'b0000000_0001101;
		Dplus[489] = 14'b0000000_0001101;
		Dplus[490] = 14'b0000000_0001101;
		Dplus[491] = 14'b0000000_0001100;
		Dplus[492] = 14'b0000000_0001100;
		Dplus[493] = 14'b0000000_0001100;
		Dplus[494] = 14'b0000000_0001100;
		Dplus[495] = 14'b0000000_0001100;
		Dplus[496] = 14'b0000000_0001100;
		Dplus[497] = 14'b0000000_0001100;
		Dplus[498] = 14'b0000000_0001100;
		Dplus[499] = 14'b0000000_0001100;
		Dplus[500] = 14'b0000000_0001100;
		Dplus[501] = 14'b0000000_0001100;
		Dplus[502] = 14'b0000000_0001100;
		Dplus[503] = 14'b0000000_0001100;
		Dplus[504] = 14'b0000000_0001100;
		Dplus[505] = 14'b0000000_0001100;
		Dplus[506] = 14'b0000000_0001100;
		Dplus[507] = 14'b0000000_0001011;
		Dplus[508] = 14'b0000000_0001011;
		Dplus[509] = 14'b0000000_0001011;
		Dplus[510] = 14'b0000000_0001011;
		Dplus[511] = 14'b0000000_0001011;
		Dplus[512] = 14'b0000000_0001011;
		Dplus[513] = 14'b0000000_0001011;
		Dplus[514] = 14'b0000000_0001011;
		Dplus[515] = 14'b0000000_0001011;
		Dplus[516] = 14'b0000000_0001011;
		Dplus[517] = 14'b0000000_0001011;
		Dplus[518] = 14'b0000000_0001011;
		Dplus[519] = 14'b0000000_0001011;
		Dplus[520] = 14'b0000000_0001011;
		Dplus[521] = 14'b0000000_0001011;
		Dplus[522] = 14'b0000000_0001011;
		Dplus[523] = 14'b0000000_0001011;
		Dplus[524] = 14'b0000000_0001011;
		Dplus[525] = 14'b0000000_0001010;
		Dplus[526] = 14'b0000000_0001010;
		Dplus[527] = 14'b0000000_0001010;
		Dplus[528] = 14'b0000000_0001010;
		Dplus[529] = 14'b0000000_0001010;
		Dplus[530] = 14'b0000000_0001010;
		Dplus[531] = 14'b0000000_0001010;
		Dplus[532] = 14'b0000000_0001010;
		Dplus[533] = 14'b0000000_0001010;
		Dplus[534] = 14'b0000000_0001010;
		Dplus[535] = 14'b0000000_0001010;
		Dplus[536] = 14'b0000000_0001010;
		Dplus[537] = 14'b0000000_0001010;
		Dplus[538] = 14'b0000000_0001010;
		Dplus[539] = 14'b0000000_0001010;
		Dplus[540] = 14'b0000000_0001010;
		Dplus[541] = 14'b0000000_0001010;
		Dplus[542] = 14'b0000000_0001010;
		Dplus[543] = 14'b0000000_0001010;
		Dplus[544] = 14'b0000000_0001001;
		Dplus[545] = 14'b0000000_0001001;
		Dplus[546] = 14'b0000000_0001001;
		Dplus[547] = 14'b0000000_0001001;
		Dplus[548] = 14'b0000000_0001001;
		Dplus[549] = 14'b0000000_0001001;
		Dplus[550] = 14'b0000000_0001001;
		Dplus[551] = 14'b0000000_0001001;
		Dplus[552] = 14'b0000000_0001001;
		Dplus[553] = 14'b0000000_0001001;
		Dplus[554] = 14'b0000000_0001001;
		Dplus[555] = 14'b0000000_0001001;
		Dplus[556] = 14'b0000000_0001001;
		Dplus[557] = 14'b0000000_0001001;
		Dplus[558] = 14'b0000000_0001001;
		Dplus[559] = 14'b0000000_0001001;
		Dplus[560] = 14'b0000000_0001001;
		Dplus[561] = 14'b0000000_0001001;
		Dplus[562] = 14'b0000000_0001001;
		Dplus[563] = 14'b0000000_0001001;
		Dplus[564] = 14'b0000000_0001001;
		Dplus[565] = 14'b0000000_0001000;
		Dplus[566] = 14'b0000000_0001000;
		Dplus[567] = 14'b0000000_0001000;
		Dplus[568] = 14'b0000000_0001000;
		Dplus[569] = 14'b0000000_0001000;
		Dplus[570] = 14'b0000000_0001000;
		Dplus[571] = 14'b0000000_0001000;
		Dplus[572] = 14'b0000000_0001000;
		Dplus[573] = 14'b0000000_0001000;
		Dplus[574] = 14'b0000000_0001000;
		Dplus[575] = 14'b0000000_0001000;
		Dplus[576] = 14'b0000000_0001000;
		Dplus[577] = 14'b0000000_0001000;
		Dplus[578] = 14'b0000000_0001000;
		Dplus[579] = 14'b0000000_0001000;
		Dplus[580] = 14'b0000000_0001000;
		Dplus[581] = 14'b0000000_0001000;
		Dplus[582] = 14'b0000000_0001000;
		Dplus[583] = 14'b0000000_0001000;
		Dplus[584] = 14'b0000000_0001000;
		Dplus[585] = 14'b0000000_0001000;
		Dplus[586] = 14'b0000000_0001000;
		Dplus[587] = 14'b0000000_0001000;
		Dplus[588] = 14'b0000000_0000111;
		Dplus[589] = 14'b0000000_0000111;
		Dplus[590] = 14'b0000000_0000111;
		Dplus[591] = 14'b0000000_0000111;
		Dplus[592] = 14'b0000000_0000111;
		Dplus[593] = 14'b0000000_0000111;
		Dplus[594] = 14'b0000000_0000111;
		Dplus[595] = 14'b0000000_0000111;
		Dplus[596] = 14'b0000000_0000111;
		Dplus[597] = 14'b0000000_0000111;
		Dplus[598] = 14'b0000000_0000111;
		Dplus[599] = 14'b0000000_0000111;
		Dplus[600] = 14'b0000000_0000111;
		Dplus[601] = 14'b0000000_0000111;
		Dplus[602] = 14'b0000000_0000111;
		Dplus[603] = 14'b0000000_0000111;
		Dplus[604] = 14'b0000000_0000111;
		Dplus[605] = 14'b0000000_0000111;
		Dplus[606] = 14'b0000000_0000111;
		Dplus[607] = 14'b0000000_0000111;
		Dplus[608] = 14'b0000000_0000111;
		Dplus[609] = 14'b0000000_0000111;
		Dplus[610] = 14'b0000000_0000111;
		Dplus[611] = 14'b0000000_0000111;
		Dplus[612] = 14'b0000000_0000111;
		Dplus[613] = 14'b0000000_0000111;
		Dplus[614] = 14'b0000000_0000111;
		Dplus[615] = 14'b0000000_0000110;
		Dplus[616] = 14'b0000000_0000110;
		Dplus[617] = 14'b0000000_0000110;
		Dplus[618] = 14'b0000000_0000110;
		Dplus[619] = 14'b0000000_0000110;
		Dplus[620] = 14'b0000000_0000110;
		Dplus[621] = 14'b0000000_0000110;
		Dplus[622] = 14'b0000000_0000110;
		Dplus[623] = 14'b0000000_0000110;
		Dplus[624] = 14'b0000000_0000110;
		Dplus[625] = 14'b0000000_0000110;
		Dplus[626] = 14'b0000000_0000110;
		Dplus[627] = 14'b0000000_0000110;
		Dplus[628] = 14'b0000000_0000110;
		Dplus[629] = 14'b0000000_0000110;
		Dplus[630] = 14'b0000000_0000110;
		Dplus[631] = 14'b0000000_0000110;
		Dplus[632] = 14'b0000000_0000110;
		Dplus[633] = 14'b0000000_0000110;
		Dplus[634] = 14'b0000000_0000110;
		Dplus[635] = 14'b0000000_0000110;
		Dplus[636] = 14'b0000000_0000110;
		Dplus[637] = 14'b0000000_0000110;
		Dplus[638] = 14'b0000000_0000110;
		Dplus[639] = 14'b0000000_0000110;
		Dplus[640] = 14'b0000000_0000110;
		Dplus[641] = 14'b0000000_0000110;
		Dplus[642] = 14'b0000000_0000110;
		Dplus[643] = 14'b0000000_0000110;
		Dplus[644] = 14'b0000000_0000110;
		Dplus[645] = 14'b0000000_0000110;
		Dplus[646] = 14'b0000000_0000110;
		Dplus[647] = 14'b0000000_0000101;
		Dplus[648] = 14'b0000000_0000101;
		Dplus[649] = 14'b0000000_0000101;
		Dplus[650] = 14'b0000000_0000101;
		Dplus[651] = 14'b0000000_0000101;
		Dplus[652] = 14'b0000000_0000101;
		Dplus[653] = 14'b0000000_0000101;
		Dplus[654] = 14'b0000000_0000101;
		Dplus[655] = 14'b0000000_0000101;
		Dplus[656] = 14'b0000000_0000101;
		Dplus[657] = 14'b0000000_0000101;
		Dplus[658] = 14'b0000000_0000101;
		Dplus[659] = 14'b0000000_0000101;
		Dplus[660] = 14'b0000000_0000101;
		Dplus[661] = 14'b0000000_0000101;
		Dplus[662] = 14'b0000000_0000101;
		Dplus[663] = 14'b0000000_0000101;
		Dplus[664] = 14'b0000000_0000101;
		Dplus[665] = 14'b0000000_0000101;
		Dplus[666] = 14'b0000000_0000101;
		Dplus[667] = 14'b0000000_0000101;
		Dplus[668] = 14'b0000000_0000101;
		Dplus[669] = 14'b0000000_0000101;
		Dplus[670] = 14'b0000000_0000101;
		Dplus[671] = 14'b0000000_0000101;
		Dplus[672] = 14'b0000000_0000101;
		Dplus[673] = 14'b0000000_0000101;
		Dplus[674] = 14'b0000000_0000101;
		Dplus[675] = 14'b0000000_0000101;
		Dplus[676] = 14'b0000000_0000101;
		Dplus[677] = 14'b0000000_0000101;
		Dplus[678] = 14'b0000000_0000101;
		Dplus[679] = 14'b0000000_0000101;
		Dplus[680] = 14'b0000000_0000101;
		Dplus[681] = 14'b0000000_0000101;
		Dplus[682] = 14'b0000000_0000101;
		Dplus[683] = 14'b0000000_0000101;
		Dplus[684] = 14'b0000000_0000100;
		Dplus[685] = 14'b0000000_0000100;
		Dplus[686] = 14'b0000000_0000100;
		Dplus[687] = 14'b0000000_0000100;
		Dplus[688] = 14'b0000000_0000100;
		Dplus[689] = 14'b0000000_0000100;
		Dplus[690] = 14'b0000000_0000100;
		Dplus[691] = 14'b0000000_0000100;
		Dplus[692] = 14'b0000000_0000100;
		Dplus[693] = 14'b0000000_0000100;
		Dplus[694] = 14'b0000000_0000100;
		Dplus[695] = 14'b0000000_0000100;
		Dplus[696] = 14'b0000000_0000100;
		Dplus[697] = 14'b0000000_0000100;
		Dplus[698] = 14'b0000000_0000100;
		Dplus[699] = 14'b0000000_0000100;
		Dplus[700] = 14'b0000000_0000100;
		Dplus[701] = 14'b0000000_0000100;
		Dplus[702] = 14'b0000000_0000100;
		Dplus[703] = 14'b0000000_0000100;
		Dplus[704] = 14'b0000000_0000100;
		Dplus[705] = 14'b0000000_0000100;
		Dplus[706] = 14'b0000000_0000100;
		Dplus[707] = 14'b0000000_0000100;
		Dplus[708] = 14'b0000000_0000100;
		Dplus[709] = 14'b0000000_0000100;
		Dplus[710] = 14'b0000000_0000100;
		Dplus[711] = 14'b0000000_0000100;
		Dplus[712] = 14'b0000000_0000100;
		Dplus[713] = 14'b0000000_0000100;
		Dplus[714] = 14'b0000000_0000100;
		Dplus[715] = 14'b0000000_0000100;
		Dplus[716] = 14'b0000000_0000100;
		Dplus[717] = 14'b0000000_0000100;
		Dplus[718] = 14'b0000000_0000100;
		Dplus[719] = 14'b0000000_0000100;
		Dplus[720] = 14'b0000000_0000100;
		Dplus[721] = 14'b0000000_0000100;
		Dplus[722] = 14'b0000000_0000100;
		Dplus[723] = 14'b0000000_0000100;
		Dplus[724] = 14'b0000000_0000100;
		Dplus[725] = 14'b0000000_0000100;
		Dplus[726] = 14'b0000000_0000100;
		Dplus[727] = 14'b0000000_0000100;
		Dplus[728] = 14'b0000000_0000100;
		Dplus[729] = 14'b0000000_0000100;
		Dplus[730] = 14'b0000000_0000100;
		Dplus[731] = 14'b0000000_0000011;
		Dplus[732] = 14'b0000000_0000011;
		Dplus[733] = 14'b0000000_0000011;
		Dplus[734] = 14'b0000000_0000011;
		Dplus[735] = 14'b0000000_0000011;
		Dplus[736] = 14'b0000000_0000011;
		Dplus[737] = 14'b0000000_0000011;
		Dplus[738] = 14'b0000000_0000011;
		Dplus[739] = 14'b0000000_0000011;
		Dplus[740] = 14'b0000000_0000011;
		Dplus[741] = 14'b0000000_0000011;
		Dplus[742] = 14'b0000000_0000011;
		Dplus[743] = 14'b0000000_0000011;
		Dplus[744] = 14'b0000000_0000011;
		Dplus[745] = 14'b0000000_0000011;
		Dplus[746] = 14'b0000000_0000011;
		Dplus[747] = 14'b0000000_0000011;
		Dplus[748] = 14'b0000000_0000011;
		Dplus[749] = 14'b0000000_0000011;
		Dplus[750] = 14'b0000000_0000011;
		Dplus[751] = 14'b0000000_0000011;
		Dplus[752] = 14'b0000000_0000011;
		Dplus[753] = 14'b0000000_0000011;
		Dplus[754] = 14'b0000000_0000011;
		Dplus[755] = 14'b0000000_0000011;
		Dplus[756] = 14'b0000000_0000011;
		Dplus[757] = 14'b0000000_0000011;
		Dplus[758] = 14'b0000000_0000011;
		Dplus[759] = 14'b0000000_0000011;
		Dplus[760] = 14'b0000000_0000011;
		Dplus[761] = 14'b0000000_0000011;
		Dplus[762] = 14'b0000000_0000011;
		Dplus[763] = 14'b0000000_0000011;
		Dplus[764] = 14'b0000000_0000011;
		Dplus[765] = 14'b0000000_0000011;
		Dplus[766] = 14'b0000000_0000011;
		Dplus[767] = 14'b0000000_0000011;
		Dplus[768] = 14'b0000000_0000011;
		Dplus[769] = 14'b0000000_0000011;
		Dplus[770] = 14'b0000000_0000011;
		Dplus[771] = 14'b0000000_0000011;
		Dplus[772] = 14'b0000000_0000011;
		Dplus[773] = 14'b0000000_0000011;
		Dplus[774] = 14'b0000000_0000011;
		Dplus[775] = 14'b0000000_0000011;
		Dplus[776] = 14'b0000000_0000011;
		Dplus[777] = 14'b0000000_0000011;
		Dplus[778] = 14'b0000000_0000011;
		Dplus[779] = 14'b0000000_0000011;
		Dplus[780] = 14'b0000000_0000011;
		Dplus[781] = 14'b0000000_0000011;
		Dplus[782] = 14'b0000000_0000011;
		Dplus[783] = 14'b0000000_0000011;
		Dplus[784] = 14'b0000000_0000011;
		Dplus[785] = 14'b0000000_0000011;
		Dplus[786] = 14'b0000000_0000011;
		Dplus[787] = 14'b0000000_0000011;
		Dplus[788] = 14'b0000000_0000011;
		Dplus[789] = 14'b0000000_0000011;
		Dplus[790] = 14'b0000000_0000011;
		Dplus[791] = 14'b0000000_0000011;
		Dplus[792] = 14'b0000000_0000011;
		Dplus[793] = 14'b0000000_0000011;
		Dplus[794] = 14'b0000000_0000010;
		Dplus[795] = 14'b0000000_0000010;
		Dplus[796] = 14'b0000000_0000010;
		Dplus[797] = 14'b0000000_0000010;
		Dplus[798] = 14'b0000000_0000010;
		Dplus[799] = 14'b0000000_0000010;
		Dplus[800] = 14'b0000000_0000010;
		Dplus[801] = 14'b0000000_0000010;
		Dplus[802] = 14'b0000000_0000010;
		Dplus[803] = 14'b0000000_0000010;
		Dplus[804] = 14'b0000000_0000010;
		Dplus[805] = 14'b0000000_0000010;
		Dplus[806] = 14'b0000000_0000010;
		Dplus[807] = 14'b0000000_0000010;
		Dplus[808] = 14'b0000000_0000010;
		Dplus[809] = 14'b0000000_0000010;
		Dplus[810] = 14'b0000000_0000010;
		Dplus[811] = 14'b0000000_0000010;
		Dplus[812] = 14'b0000000_0000010;
		Dplus[813] = 14'b0000000_0000010;
		Dplus[814] = 14'b0000000_0000010;
		Dplus[815] = 14'b0000000_0000010;
		Dplus[816] = 14'b0000000_0000010;
		Dplus[817] = 14'b0000000_0000010;
		Dplus[818] = 14'b0000000_0000010;
		Dplus[819] = 14'b0000000_0000010;
		Dplus[820] = 14'b0000000_0000010;
		Dplus[821] = 14'b0000000_0000010;
		Dplus[822] = 14'b0000000_0000010;
		Dplus[823] = 14'b0000000_0000010;
		Dplus[824] = 14'b0000000_0000010;
		Dplus[825] = 14'b0000000_0000010;
		Dplus[826] = 14'b0000000_0000010;
		Dplus[827] = 14'b0000000_0000010;
		Dplus[828] = 14'b0000000_0000010;
		Dplus[829] = 14'b0000000_0000010;
		Dplus[830] = 14'b0000000_0000010;
		Dplus[831] = 14'b0000000_0000010;
		Dplus[832] = 14'b0000000_0000010;
		Dplus[833] = 14'b0000000_0000010;
		Dplus[834] = 14'b0000000_0000010;
		Dplus[835] = 14'b0000000_0000010;
		Dplus[836] = 14'b0000000_0000010;
		Dplus[837] = 14'b0000000_0000010;
		Dplus[838] = 14'b0000000_0000010;
		Dplus[839] = 14'b0000000_0000010;
		Dplus[840] = 14'b0000000_0000010;
		Dplus[841] = 14'b0000000_0000010;
		Dplus[842] = 14'b0000000_0000010;
		Dplus[843] = 14'b0000000_0000010;
		Dplus[844] = 14'b0000000_0000010;
		Dplus[845] = 14'b0000000_0000010;
		Dplus[846] = 14'b0000000_0000010;
		Dplus[847] = 14'b0000000_0000010;
		Dplus[848] = 14'b0000000_0000010;
		Dplus[849] = 14'b0000000_0000010;
		Dplus[850] = 14'b0000000_0000010;
		Dplus[851] = 14'b0000000_0000010;
		Dplus[852] = 14'b0000000_0000010;
		Dplus[853] = 14'b0000000_0000010;
		Dplus[854] = 14'b0000000_0000010;
		Dplus[855] = 14'b0000000_0000010;
		Dplus[856] = 14'b0000000_0000010;
		Dplus[857] = 14'b0000000_0000010;
		Dplus[858] = 14'b0000000_0000010;
		Dplus[859] = 14'b0000000_0000010;
		Dplus[860] = 14'b0000000_0000010;
		Dplus[861] = 14'b0000000_0000010;
		Dplus[862] = 14'b0000000_0000010;
		Dplus[863] = 14'b0000000_0000010;
		Dplus[864] = 14'b0000000_0000010;
		Dplus[865] = 14'b0000000_0000010;
		Dplus[866] = 14'b0000000_0000010;
		Dplus[867] = 14'b0000000_0000010;
		Dplus[868] = 14'b0000000_0000010;
		Dplus[869] = 14'b0000000_0000010;
		Dplus[870] = 14'b0000000_0000010;
		Dplus[871] = 14'b0000000_0000010;
		Dplus[872] = 14'b0000000_0000010;
		Dplus[873] = 14'b0000000_0000010;
		Dplus[874] = 14'b0000000_0000010;
		Dplus[875] = 14'b0000000_0000010;
		Dplus[876] = 14'b0000000_0000010;
		Dplus[877] = 14'b0000000_0000010;
		Dplus[878] = 14'b0000000_0000010;
		Dplus[879] = 14'b0000000_0000010;
		Dplus[880] = 14'b0000000_0000010;
		Dplus[881] = 14'b0000000_0000010;
		Dplus[882] = 14'b0000000_0000010;
		Dplus[883] = 14'b0000000_0000010;
		Dplus[884] = 14'b0000000_0000010;
		Dplus[885] = 14'b0000000_0000010;
		Dplus[886] = 14'b0000000_0000010;
		Dplus[887] = 14'b0000000_0000010;
		Dplus[888] = 14'b0000000_0000010;
		Dplus[889] = 14'b0000000_0000001;
		Dplus[890] = 14'b0000000_0000001;
		Dplus[891] = 14'b0000000_0000001;
		Dplus[892] = 14'b0000000_0000001;
		Dplus[893] = 14'b0000000_0000001;
		Dplus[894] = 14'b0000000_0000001;
		Dplus[895] = 14'b0000000_0000001;
		Dplus[896] = 14'b0000000_0000001;
		Dplus[897] = 14'b0000000_0000001;
		Dplus[898] = 14'b0000000_0000001;
		Dplus[899] = 14'b0000000_0000001;
		Dplus[900] = 14'b0000000_0000001;
		Dplus[901] = 14'b0000000_0000001;
		Dplus[902] = 14'b0000000_0000001;
		Dplus[903] = 14'b0000000_0000001;
		Dplus[904] = 14'b0000000_0000001;
		Dplus[905] = 14'b0000000_0000001;
		Dplus[906] = 14'b0000000_0000001;
		Dplus[907] = 14'b0000000_0000001;
		Dplus[908] = 14'b0000000_0000001;
		Dplus[909] = 14'b0000000_0000001;
		Dplus[910] = 14'b0000000_0000001;
		Dplus[911] = 14'b0000000_0000001;
		Dplus[912] = 14'b0000000_0000001;
		Dplus[913] = 14'b0000000_0000001;
		Dplus[914] = 14'b0000000_0000001;
		Dplus[915] = 14'b0000000_0000001;
		Dplus[916] = 14'b0000000_0000001;
		Dplus[917] = 14'b0000000_0000001;
		Dplus[918] = 14'b0000000_0000001;
		Dplus[919] = 14'b0000000_0000001;
		Dplus[920] = 14'b0000000_0000001;
		Dplus[921] = 14'b0000000_0000001;
		Dplus[922] = 14'b0000000_0000001;
		Dplus[923] = 14'b0000000_0000001;
		Dplus[924] = 14'b0000000_0000001;
		Dplus[925] = 14'b0000000_0000001;
		Dplus[926] = 14'b0000000_0000001;
		Dplus[927] = 14'b0000000_0000001;
		Dplus[928] = 14'b0000000_0000001;
		Dplus[929] = 14'b0000000_0000001;
		Dplus[930] = 14'b0000000_0000001;
		Dplus[931] = 14'b0000000_0000001;
		Dplus[932] = 14'b0000000_0000001;
		Dplus[933] = 14'b0000000_0000001;
		Dplus[934] = 14'b0000000_0000001;
		Dplus[935] = 14'b0000000_0000001;
		Dplus[936] = 14'b0000000_0000001;
		Dplus[937] = 14'b0000000_0000001;
		Dplus[938] = 14'b0000000_0000001;
		Dplus[939] = 14'b0000000_0000001;
		Dplus[940] = 14'b0000000_0000001;
		Dplus[941] = 14'b0000000_0000001;
		Dplus[942] = 14'b0000000_0000001;
		Dplus[943] = 14'b0000000_0000001;
		Dplus[944] = 14'b0000000_0000001;
		Dplus[945] = 14'b0000000_0000001;
		Dplus[946] = 14'b0000000_0000001;
		Dplus[947] = 14'b0000000_0000001;
		Dplus[948] = 14'b0000000_0000001;
		Dplus[949] = 14'b0000000_0000001;
		Dplus[950] = 14'b0000000_0000001;
		Dplus[951] = 14'b0000000_0000001;
		Dplus[952] = 14'b0000000_0000001;
		Dplus[953] = 14'b0000000_0000001;
		Dplus[954] = 14'b0000000_0000001;
		Dplus[955] = 14'b0000000_0000001;
		Dplus[956] = 14'b0000000_0000001;
		Dplus[957] = 14'b0000000_0000001;
		Dplus[958] = 14'b0000000_0000001;
		Dplus[959] = 14'b0000000_0000001;
		Dplus[960] = 14'b0000000_0000001;
		Dplus[961] = 14'b0000000_0000001;
		Dplus[962] = 14'b0000000_0000001;
		Dplus[963] = 14'b0000000_0000001;
		Dplus[964] = 14'b0000000_0000001;
		Dplus[965] = 14'b0000000_0000001;
		Dplus[966] = 14'b0000000_0000001;
		Dplus[967] = 14'b0000000_0000001;
		Dplus[968] = 14'b0000000_0000001;
		Dplus[969] = 14'b0000000_0000001;
		Dplus[970] = 14'b0000000_0000001;
		Dplus[971] = 14'b0000000_0000001;
		Dplus[972] = 14'b0000000_0000001;
		Dplus[973] = 14'b0000000_0000001;
		Dplus[974] = 14'b0000000_0000001;
		Dplus[975] = 14'b0000000_0000001;
		Dplus[976] = 14'b0000000_0000001;
		Dplus[977] = 14'b0000000_0000001;
		Dplus[978] = 14'b0000000_0000001;
		Dplus[979] = 14'b0000000_0000001;
		Dplus[980] = 14'b0000000_0000001;
		Dplus[981] = 14'b0000000_0000001;
		Dplus[982] = 14'b0000000_0000001;
		Dplus[983] = 14'b0000000_0000001;
		Dplus[984] = 14'b0000000_0000001;
		Dplus[985] = 14'b0000000_0000001;
		Dplus[986] = 14'b0000000_0000001;
		Dplus[987] = 14'b0000000_0000001;
		Dplus[988] = 14'b0000000_0000001;
		Dplus[989] = 14'b0000000_0000001;
		Dplus[990] = 14'b0000000_0000001;
		Dplus[991] = 14'b0000000_0000001;
		Dplus[992] = 14'b0000000_0000001;
		Dplus[993] = 14'b0000000_0000001;
		Dplus[994] = 14'b0000000_0000001;
		Dplus[995] = 14'b0000000_0000001;
		Dplus[996] = 14'b0000000_0000001;
		Dplus[997] = 14'b0000000_0000001;
		Dplus[998] = 14'b0000000_0000001;
		Dplus[999] = 14'b0000000_0000001;
		Dplus[1000] = 14'b0000000_0000001;
		Dplus[1001] = 14'b0000000_0000001;
		Dplus[1002] = 14'b0000000_0000001;
		Dplus[1003] = 14'b0000000_0000001;
		Dplus[1004] = 14'b0000000_0000001;
		Dplus[1005] = 14'b0000000_0000001;
		Dplus[1006] = 14'b0000000_0000001;
		Dplus[1007] = 14'b0000000_0000001;
		Dplus[1008] = 14'b0000000_0000001;
		Dplus[1009] = 14'b0000000_0000001;
		Dplus[1010] = 14'b0000000_0000001;
		Dplus[1011] = 14'b0000000_0000001;
		Dplus[1012] = 14'b0000000_0000001;
		Dplus[1013] = 14'b0000000_0000001;
		Dplus[1014] = 14'b0000000_0000001;
		Dplus[1015] = 14'b0000000_0000001;
		Dplus[1016] = 14'b0000000_0000001;
		Dplus[1017] = 14'b0000000_0000001;
		Dplus[1018] = 14'b0000000_0000001;
		Dplus[1019] = 14'b0000000_0000001;
		Dplus[1020] = 14'b0000000_0000001;
		Dplus[1021] = 14'b0000000_0000001;
		Dplus[1022] = 14'b0000000_0000001;
		Dplus[1023] = 14'b0000000_0000001;
		Dplus[1024] = 14'b0000000_0000001;
		Dplus[1025] = 14'b0000000_0000001;
		Dplus[1026] = 14'b0000000_0000001;
		Dplus[1027] = 14'b0000000_0000001;
		Dplus[1028] = 14'b0000000_0000001;
		Dplus[1029] = 14'b0000000_0000001;
		Dplus[1030] = 14'b0000000_0000001;
		Dplus[1031] = 14'b0000000_0000001;
		Dplus[1032] = 14'b0000000_0000001;
		Dplus[1033] = 14'b0000000_0000001;
		Dplus[1034] = 14'b0000000_0000001;
		Dplus[1035] = 14'b0000000_0000001;
		Dplus[1036] = 14'b0000000_0000001;
		Dplus[1037] = 14'b0000000_0000001;
		Dplus[1038] = 14'b0000000_0000001;
		Dplus[1039] = 14'b0000000_0000001;
		Dplus[1040] = 14'b0000000_0000001;
		Dplus[1041] = 14'b0000000_0000001;
		Dplus[1042] = 14'b0000000_0000001;
		Dplus[1043] = 14'b0000000_0000001;
		Dplus[1044] = 14'b0000000_0000001;
		Dplus[1045] = 14'b0000000_0000001;
		Dplus[1046] = 14'b0000000_0000001;
		Dplus[1047] = 14'b0000000_0000001;
		Dplus[1048] = 14'b0000000_0000001;
		Dplus[1049] = 14'b0000000_0000001;
		Dplus[1050] = 14'b0000000_0000001;
		Dplus[1051] = 14'b0000000_0000001;
		Dplus[1052] = 14'b0000000_0000001;
		Dplus[1053] = 14'b0000000_0000001;
		Dplus[1054] = 14'b0000000_0000001;
		Dplus[1055] = 14'b0000000_0000001;
		Dplus[1056] = 14'b0000000_0000001;
		Dplus[1057] = 14'b0000000_0000001;
		Dplus[1058] = 14'b0000000_0000001;
		Dplus[1059] = 14'b0000000_0000001;
		Dplus[1060] = 14'b0000000_0000001;
		Dplus[1061] = 14'b0000000_0000001;
		Dplus[1062] = 14'b0000000_0000001;
		Dplus[1063] = 14'b0000000_0000001;
		Dplus[1064] = 14'b0000000_0000001;
		Dplus[1065] = 14'b0000000_0000001;
		Dplus[1066] = 14'b0000000_0000001;
		Dplus[1067] = 14'b0000000_0000001;
		Dplus[1068] = 14'b0000000_0000001;
		Dplus[1069] = 14'b0000000_0000001;
		Dplus[1070] = 14'b0000000_0000001;
		Dplus[1071] = 14'b0000000_0000001;
		Dplus[1072] = 14'b0000000_0000001;
		Dplus[1073] = 14'b0000000_0000001;
		Dplus[1074] = 14'b0000000_0000001;
		Dplus[1075] = 14'b0000000_0000001;
		Dplus[1076] = 14'b0000000_0000001;
		Dplus[1077] = 14'b0000000_0000001;
		Dplus[1078] = 14'b0000000_0000001;
		Dplus[1079] = 14'b0000000_0000001;
		Dplus[1080] = 14'b0000000_0000001;
		Dplus[1081] = 14'b0000000_0000001;
		Dplus[1082] = 14'b0000000_0000001;
		Dplus[1083] = 14'b0000000_0000001;
		Dplus[1084] = 14'b0000000_0000001;
		Dplus[1085] = 14'b0000000_0000001;
		Dplus[1086] = 14'b0000000_0000001;
		Dplus[1087] = 14'b0000000_0000001;
		Dplus[1088] = 14'b0000000_0000001;
		Dplus[1089] = 14'b0000000_0000001;
		Dplus[1090] = 14'b0000000_0000001;
		Dplus[1091] = 14'b0000000_0000001;
		Dplus[1092] = 14'b0000000_0000000;
		Dplus[1093] = 14'b0000000_0000000;
		Dplus[1094] = 14'b0000000_0000000;
		Dplus[1095] = 14'b0000000_0000000;
		Dplus[1096] = 14'b0000000_0000000;
		Dplus[1097] = 14'b0000000_0000000;
		Dplus[1098] = 14'b0000000_0000000;
		Dplus[1099] = 14'b0000000_0000000;
		Dplus[1100] = 14'b0000000_0000000;
		Dplus[1101] = 14'b0000000_0000000;
		Dplus[1102] = 14'b0000000_0000000;
		Dplus[1103] = 14'b0000000_0000000;
		Dplus[1104] = 14'b0000000_0000000;
		Dplus[1105] = 14'b0000000_0000000;
		Dplus[1106] = 14'b0000000_0000000;
		Dplus[1107] = 14'b0000000_0000000;
		Dplus[1108] = 14'b0000000_0000000;
		Dplus[1109] = 14'b0000000_0000000;
		Dplus[1110] = 14'b0000000_0000000;
		Dplus[1111] = 14'b0000000_0000000;
		Dplus[1112] = 14'b0000000_0000000;
		Dplus[1113] = 14'b0000000_0000000;
		Dplus[1114] = 14'b0000000_0000000;
		Dplus[1115] = 14'b0000000_0000000;
		Dplus[1116] = 14'b0000000_0000000;
		Dplus[1117] = 14'b0000000_0000000;
		Dplus[1118] = 14'b0000000_0000000;
		Dplus[1119] = 14'b0000000_0000000;
		Dplus[1120] = 14'b0000000_0000000;
		Dplus[1121] = 14'b0000000_0000000;
		Dplus[1122] = 14'b0000000_0000000;
		Dplus[1123] = 14'b0000000_0000000;
		Dplus[1124] = 14'b0000000_0000000;
		Dplus[1125] = 14'b0000000_0000000;
		Dplus[1126] = 14'b0000000_0000000;
		Dplus[1127] = 14'b0000000_0000000;
		Dplus[1128] = 14'b0000000_0000000;
		Dplus[1129] = 14'b0000000_0000000;
		Dplus[1130] = 14'b0000000_0000000;
		Dplus[1131] = 14'b0000000_0000000;
		Dplus[1132] = 14'b0000000_0000000;
		Dplus[1133] = 14'b0000000_0000000;
		Dplus[1134] = 14'b0000000_0000000;
		Dplus[1135] = 14'b0000000_0000000;
		Dplus[1136] = 14'b0000000_0000000;
		Dplus[1137] = 14'b0000000_0000000;
		Dplus[1138] = 14'b0000000_0000000;
		Dplus[1139] = 14'b0000000_0000000;
		Dplus[1140] = 14'b0000000_0000000;
		Dplus[1141] = 14'b0000000_0000000;
		Dplus[1142] = 14'b0000000_0000000;
		Dplus[1143] = 14'b0000000_0000000;
		Dplus[1144] = 14'b0000000_0000000;
		Dplus[1145] = 14'b0000000_0000000;
		Dplus[1146] = 14'b0000000_0000000;
		Dplus[1147] = 14'b0000000_0000000;
		Dplus[1148] = 14'b0000000_0000000;
		Dplus[1149] = 14'b0000000_0000000;
		Dplus[1150] = 14'b0000000_0000000;
		Dplus[1151] = 14'b0000000_0000000;
		Dplus[1152] = 14'b0000000_0000000;
		Dplus[1153] = 14'b0000000_0000000;
		Dplus[1154] = 14'b0000000_0000000;
		Dplus[1155] = 14'b0000000_0000000;
		Dplus[1156] = 14'b0000000_0000000;
		Dplus[1157] = 14'b0000000_0000000;
		Dplus[1158] = 14'b0000000_0000000;
		Dplus[1159] = 14'b0000000_0000000;
		Dplus[1160] = 14'b0000000_0000000;
		Dplus[1161] = 14'b0000000_0000000;
		Dplus[1162] = 14'b0000000_0000000;
		Dplus[1163] = 14'b0000000_0000000;
		Dplus[1164] = 14'b0000000_0000000;
		Dplus[1165] = 14'b0000000_0000000;
		Dplus[1166] = 14'b0000000_0000000;
		Dplus[1167] = 14'b0000000_0000000;
		Dplus[1168] = 14'b0000000_0000000;
		Dplus[1169] = 14'b0000000_0000000;
		Dplus[1170] = 14'b0000000_0000000;
		Dplus[1171] = 14'b0000000_0000000;
		Dplus[1172] = 14'b0000000_0000000;
		Dplus[1173] = 14'b0000000_0000000;
		Dplus[1174] = 14'b0000000_0000000;
		Dplus[1175] = 14'b0000000_0000000;
		Dplus[1176] = 14'b0000000_0000000;
		Dplus[1177] = 14'b0000000_0000000;
		Dplus[1178] = 14'b0000000_0000000;
		Dplus[1179] = 14'b0000000_0000000;
		Dplus[1180] = 14'b0000000_0000000;
		Dplus[1181] = 14'b0000000_0000000;
		Dplus[1182] = 14'b0000000_0000000;
		Dplus[1183] = 14'b0000000_0000000;
		Dplus[1184] = 14'b0000000_0000000;
		Dplus[1185] = 14'b0000000_0000000;
		Dplus[1186] = 14'b0000000_0000000;
		Dplus[1187] = 14'b0000000_0000000;
		Dplus[1188] = 14'b0000000_0000000;
		Dplus[1189] = 14'b0000000_0000000;
		Dplus[1190] = 14'b0000000_0000000;
		Dplus[1191] = 14'b0000000_0000000;
		Dplus[1192] = 14'b0000000_0000000;
		Dplus[1193] = 14'b0000000_0000000;
		Dplus[1194] = 14'b0000000_0000000;
		Dplus[1195] = 14'b0000000_0000000;
		Dplus[1196] = 14'b0000000_0000000;
		Dplus[1197] = 14'b0000000_0000000;
		Dplus[1198] = 14'b0000000_0000000;
		Dplus[1199] = 14'b0000000_0000000;
		Dplus[1200] = 14'b0000000_0000000;
		Dplus[1201] = 14'b0000000_0000000;
		Dplus[1202] = 14'b0000000_0000000;
		Dplus[1203] = 14'b0000000_0000000;
		Dplus[1204] = 14'b0000000_0000000;
		Dplus[1205] = 14'b0000000_0000000;
		Dplus[1206] = 14'b0000000_0000000;
		Dplus[1207] = 14'b0000000_0000000;
		Dplus[1208] = 14'b0000000_0000000;
		Dplus[1209] = 14'b0000000_0000000;
		Dplus[1210] = 14'b0000000_0000000;
		Dplus[1211] = 14'b0000000_0000000;
		Dplus[1212] = 14'b0000000_0000000;
		Dplus[1213] = 14'b0000000_0000000;
		Dplus[1214] = 14'b0000000_0000000;
		Dplus[1215] = 14'b0000000_0000000;
		Dplus[1216] = 14'b0000000_0000000;
		Dplus[1217] = 14'b0000000_0000000;
		Dplus[1218] = 14'b0000000_0000000;
		Dplus[1219] = 14'b0000000_0000000;
		Dplus[1220] = 14'b0000000_0000000;
		Dplus[1221] = 14'b0000000_0000000;
		Dplus[1222] = 14'b0000000_0000000;
		Dplus[1223] = 14'b0000000_0000000;
		Dplus[1224] = 14'b0000000_0000000;
		Dplus[1225] = 14'b0000000_0000000;
		Dplus[1226] = 14'b0000000_0000000;
		Dplus[1227] = 14'b0000000_0000000;
		Dplus[1228] = 14'b0000000_0000000;
		Dplus[1229] = 14'b0000000_0000000;
		Dplus[1230] = 14'b0000000_0000000;
		Dplus[1231] = 14'b0000000_0000000;
		Dplus[1232] = 14'b0000000_0000000;
		Dplus[1233] = 14'b0000000_0000000;
		Dplus[1234] = 14'b0000000_0000000;
		Dplus[1235] = 14'b0000000_0000000;
		Dplus[1236] = 14'b0000000_0000000;
		Dplus[1237] = 14'b0000000_0000000;
		Dplus[1238] = 14'b0000000_0000000;
		Dplus[1239] = 14'b0000000_0000000;
		Dplus[1240] = 14'b0000000_0000000;
		Dplus[1241] = 14'b0000000_0000000;
		Dplus[1242] = 14'b0000000_0000000;
		Dplus[1243] = 14'b0000000_0000000;
		Dplus[1244] = 14'b0000000_0000000;
		Dplus[1245] = 14'b0000000_0000000;
		Dplus[1246] = 14'b0000000_0000000;
		Dplus[1247] = 14'b0000000_0000000;
		Dplus[1248] = 14'b0000000_0000000;
		Dplus[1249] = 14'b0000000_0000000;
		Dplus[1250] = 14'b0000000_0000000;
		Dplus[1251] = 14'b0000000_0000000;
		Dplus[1252] = 14'b0000000_0000000;
		Dplus[1253] = 14'b0000000_0000000;
		Dplus[1254] = 14'b0000000_0000000;
		Dplus[1255] = 14'b0000000_0000000;
		Dplus[1256] = 14'b0000000_0000000;
		Dplus[1257] = 14'b0000000_0000000;
		Dplus[1258] = 14'b0000000_0000000;
		Dplus[1259] = 14'b0000000_0000000;
		Dplus[1260] = 14'b0000000_0000000;
		Dplus[1261] = 14'b0000000_0000000;
		Dplus[1262] = 14'b0000000_0000000;
		Dplus[1263] = 14'b0000000_0000000;
		Dplus[1264] = 14'b0000000_0000000;
		Dplus[1265] = 14'b0000000_0000000;
		Dplus[1266] = 14'b0000000_0000000;
		Dplus[1267] = 14'b0000000_0000000;
		Dplus[1268] = 14'b0000000_0000000;
		Dplus[1269] = 14'b0000000_0000000;
		Dplus[1270] = 14'b0000000_0000000;
		Dplus[1271] = 14'b0000000_0000000;
		Dplus[1272] = 14'b0000000_0000000;
		Dplus[1273] = 14'b0000000_0000000;
		Dplus[1274] = 14'b0000000_0000000;
		Dplus[1275] = 14'b0000000_0000000;
		Dplus[1276] = 14'b0000000_0000000;
		Dplus[1277] = 14'b0000000_0000000;
		Dplus[1278] = 14'b0000000_0000000;
		Dplus[1279] = 14'b0000000_0000000;
		Dplus[1280] = 14'b0000000_0000000;
		Dplus[1281] = 14'b0000000_0000000;
		Dplus[1282] = 14'b0000000_0000000;
		Dplus[1283] = 14'b0000000_0000000;
		Dplus[1284] = 14'b0000000_0000000;
		Dplus[1285] = 14'b0000000_0000000;
		Dplus[1286] = 14'b0000000_0000000;
		Dplus[1287] = 14'b0000000_0000000;
		Dplus[1288] = 14'b0000000_0000000;
		Dplus[1289] = 14'b0000000_0000000;
		Dplus[1290] = 14'b0000000_0000000;
		Dplus[1291] = 14'b0000000_0000000;
		Dplus[1292] = 14'b0000000_0000000;
		Dplus[1293] = 14'b0000000_0000000;
		Dplus[1294] = 14'b0000000_0000000;
		Dplus[1295] = 14'b0000000_0000000;
		Dplus[1296] = 14'b0000000_0000000;
		Dplus[1297] = 14'b0000000_0000000;
		Dplus[1298] = 14'b0000000_0000000;
		Dplus[1299] = 14'b0000000_0000000;
		Dplus[1300] = 14'b0000000_0000000;
		Dplus[1301] = 14'b0000000_0000000;
		Dplus[1302] = 14'b0000000_0000000;
		Dplus[1303] = 14'b0000000_0000000;
		Dplus[1304] = 14'b0000000_0000000;
		Dplus[1305] = 14'b0000000_0000000;
		Dplus[1306] = 14'b0000000_0000000;
		Dplus[1307] = 14'b0000000_0000000;
		Dplus[1308] = 14'b0000000_0000000;
		Dplus[1309] = 14'b0000000_0000000;
		Dplus[1310] = 14'b0000000_0000000;
		Dplus[1311] = 14'b0000000_0000000;
		Dplus[1312] = 14'b0000000_0000000;
		Dplus[1313] = 14'b0000000_0000000;
		Dplus[1314] = 14'b0000000_0000000;
		Dplus[1315] = 14'b0000000_0000000;
		Dplus[1316] = 14'b0000000_0000000;
		Dplus[1317] = 14'b0000000_0000000;
		Dplus[1318] = 14'b0000000_0000000;
		Dplus[1319] = 14'b0000000_0000000;
		Dplus[1320] = 14'b0000000_0000000;
		Dplus[1321] = 14'b0000000_0000000;
		Dplus[1322] = 14'b0000000_0000000;
		Dplus[1323] = 14'b0000000_0000000;
		Dplus[1324] = 14'b0000000_0000000;
		Dplus[1325] = 14'b0000000_0000000;
		Dplus[1326] = 14'b0000000_0000000;
		Dplus[1327] = 14'b0000000_0000000;
		Dplus[1328] = 14'b0000000_0000000;
		Dplus[1329] = 14'b0000000_0000000;
		Dplus[1330] = 14'b0000000_0000000;
		Dplus[1331] = 14'b0000000_0000000;
		Dplus[1332] = 14'b0000000_0000000;
		Dplus[1333] = 14'b0000000_0000000;
		Dplus[1334] = 14'b0000000_0000000;
		Dplus[1335] = 14'b0000000_0000000;
		Dplus[1336] = 14'b0000000_0000000;
		Dplus[1337] = 14'b0000000_0000000;
		Dplus[1338] = 14'b0000000_0000000;
		Dplus[1339] = 14'b0000000_0000000;
		Dplus[1340] = 14'b0000000_0000000;
		Dplus[1341] = 14'b0000000_0000000;
		Dplus[1342] = 14'b0000000_0000000;
		Dplus[1343] = 14'b0000000_0000000;
		Dplus[1344] = 14'b0000000_0000000;
		Dplus[1345] = 14'b0000000_0000000;
		Dplus[1346] = 14'b0000000_0000000;
		Dplus[1347] = 14'b0000000_0000000;
		Dplus[1348] = 14'b0000000_0000000;
		Dplus[1349] = 14'b0000000_0000000;
		Dplus[1350] = 14'b0000000_0000000;
		Dplus[1351] = 14'b0000000_0000000;
		Dplus[1352] = 14'b0000000_0000000;
		Dplus[1353] = 14'b0000000_0000000;
		Dplus[1354] = 14'b0000000_0000000;
		Dplus[1355] = 14'b0000000_0000000;
		Dplus[1356] = 14'b0000000_0000000;
		Dplus[1357] = 14'b0000000_0000000;
		Dplus[1358] = 14'b0000000_0000000;
		Dplus[1359] = 14'b0000000_0000000;
		Dplus[1360] = 14'b0000000_0000000;
		Dplus[1361] = 14'b0000000_0000000;
		Dplus[1362] = 14'b0000000_0000000;
		Dplus[1363] = 14'b0000000_0000000;
		Dplus[1364] = 14'b0000000_0000000;
		Dplus[1365] = 14'b0000000_0000000;
		Dplus[1366] = 14'b0000000_0000000;
		Dplus[1367] = 14'b0000000_0000000;
		Dplus[1368] = 14'b0000000_0000000;
		Dplus[1369] = 14'b0000000_0000000;
		Dplus[1370] = 14'b0000000_0000000;
		Dplus[1371] = 14'b0000000_0000000;
		Dplus[1372] = 14'b0000000_0000000;
		Dplus[1373] = 14'b0000000_0000000;
		Dplus[1374] = 14'b0000000_0000000;
		Dplus[1375] = 14'b0000000_0000000;
		Dplus[1376] = 14'b0000000_0000000;
		Dplus[1377] = 14'b0000000_0000000;
		Dplus[1378] = 14'b0000000_0000000;
		Dplus[1379] = 14'b0000000_0000000;
		Dplus[1380] = 14'b0000000_0000000;
		Dplus[1381] = 14'b0000000_0000000;
		Dplus[1382] = 14'b0000000_0000000;
		Dplus[1383] = 14'b0000000_0000000;
		Dplus[1384] = 14'b0000000_0000000;
		Dplus[1385] = 14'b0000000_0000000;
		Dplus[1386] = 14'b0000000_0000000;
		Dplus[1387] = 14'b0000000_0000000;
		Dplus[1388] = 14'b0000000_0000000;
		Dplus[1389] = 14'b0000000_0000000;
		Dplus[1390] = 14'b0000000_0000000;
		Dplus[1391] = 14'b0000000_0000000;
		Dplus[1392] = 14'b0000000_0000000;
		Dplus[1393] = 14'b0000000_0000000;
		Dplus[1394] = 14'b0000000_0000000;
		Dplus[1395] = 14'b0000000_0000000;
		Dplus[1396] = 14'b0000000_0000000;
		Dplus[1397] = 14'b0000000_0000000;
		Dplus[1398] = 14'b0000000_0000000;
		Dplus[1399] = 14'b0000000_0000000;
		Dplus[1400] = 14'b0000000_0000000;
		Dplus[1401] = 14'b0000000_0000000;
		Dplus[1402] = 14'b0000000_0000000;
		Dplus[1403] = 14'b0000000_0000000;
		Dplus[1404] = 14'b0000000_0000000;
		Dplus[1405] = 14'b0000000_0000000;
		Dplus[1406] = 14'b0000000_0000000;
		Dplus[1407] = 14'b0000000_0000000;
		Dplus[1408] = 14'b0000000_0000000;
		Dplus[1409] = 14'b0000000_0000000;
		Dplus[1410] = 14'b0000000_0000000;
		Dplus[1411] = 14'b0000000_0000000;
		Dplus[1412] = 14'b0000000_0000000;
		Dplus[1413] = 14'b0000000_0000000;
		Dplus[1414] = 14'b0000000_0000000;
		Dplus[1415] = 14'b0000000_0000000;
		Dplus[1416] = 14'b0000000_0000000;
		Dplus[1417] = 14'b0000000_0000000;
		Dplus[1418] = 14'b0000000_0000000;
		Dplus[1419] = 14'b0000000_0000000;
		Dplus[1420] = 14'b0000000_0000000;
		Dplus[1421] = 14'b0000000_0000000;
		Dplus[1422] = 14'b0000000_0000000;
		Dplus[1423] = 14'b0000000_0000000;
		Dplus[1424] = 14'b0000000_0000000;
		Dplus[1425] = 14'b0000000_0000000;
		Dplus[1426] = 14'b0000000_0000000;
		Dplus[1427] = 14'b0000000_0000000;
		Dplus[1428] = 14'b0000000_0000000;
		Dplus[1429] = 14'b0000000_0000000;
		Dplus[1430] = 14'b0000000_0000000;
		Dplus[1431] = 14'b0000000_0000000;
		Dplus[1432] = 14'b0000000_0000000;
		Dplus[1433] = 14'b0000000_0000000;
		Dplus[1434] = 14'b0000000_0000000;
		Dplus[1435] = 14'b0000000_0000000;
		Dplus[1436] = 14'b0000000_0000000;
		Dplus[1437] = 14'b0000000_0000000;
		Dplus[1438] = 14'b0000000_0000000;
		Dplus[1439] = 14'b0000000_0000000;
		Dplus[1440] = 14'b0000000_0000000;
		Dplus[1441] = 14'b0000000_0000000;
		Dplus[1442] = 14'b0000000_0000000;
		Dplus[1443] = 14'b0000000_0000000;
		Dplus[1444] = 14'b0000000_0000000;
		Dplus[1445] = 14'b0000000_0000000;
		Dplus[1446] = 14'b0000000_0000000;
		Dplus[1447] = 14'b0000000_0000000;
		Dplus[1448] = 14'b0000000_0000000;
		Dplus[1449] = 14'b0000000_0000000;
		Dplus[1450] = 14'b0000000_0000000;
		Dplus[1451] = 14'b0000000_0000000;
		Dplus[1452] = 14'b0000000_0000000;
		Dplus[1453] = 14'b0000000_0000000;
		Dplus[1454] = 14'b0000000_0000000;
		Dplus[1455] = 14'b0000000_0000000;
		Dplus[1456] = 14'b0000000_0000000;
		Dplus[1457] = 14'b0000000_0000000;
		Dplus[1458] = 14'b0000000_0000000;
		Dplus[1459] = 14'b0000000_0000000;
		Dplus[1460] = 14'b0000000_0000000;
		Dplus[1461] = 14'b0000000_0000000;
		Dplus[1462] = 14'b0000000_0000000;
		Dplus[1463] = 14'b0000000_0000000;
		Dplus[1464] = 14'b0000000_0000000;
		Dplus[1465] = 14'b0000000_0000000;
		Dplus[1466] = 14'b0000000_0000000;
		Dplus[1467] = 14'b0000000_0000000;
		Dplus[1468] = 14'b0000000_0000000;
		Dplus[1469] = 14'b0000000_0000000;
		Dplus[1470] = 14'b0000000_0000000;
		Dplus[1471] = 14'b0000000_0000000;
		Dplus[1472] = 14'b0000000_0000000;
		Dplus[1473] = 14'b0000000_0000000;
		Dplus[1474] = 14'b0000000_0000000;
		Dplus[1475] = 14'b0000000_0000000;
		Dplus[1476] = 14'b0000000_0000000;
		Dplus[1477] = 14'b0000000_0000000;
		Dplus[1478] = 14'b0000000_0000000;
		Dplus[1479] = 14'b0000000_0000000;
		Dplus[1480] = 14'b0000000_0000000;
		Dplus[1481] = 14'b0000000_0000000;
		Dplus[1482] = 14'b0000000_0000000;
		Dplus[1483] = 14'b0000000_0000000;
		Dplus[1484] = 14'b0000000_0000000;
		Dplus[1485] = 14'b0000000_0000000;
		Dplus[1486] = 14'b0000000_0000000;
		Dplus[1487] = 14'b0000000_0000000;
		Dplus[1488] = 14'b0000000_0000000;
		Dplus[1489] = 14'b0000000_0000000;
		Dplus[1490] = 14'b0000000_0000000;
		Dplus[1491] = 14'b0000000_0000000;
		Dplus[1492] = 14'b0000000_0000000;
		Dplus[1493] = 14'b0000000_0000000;
		Dplus[1494] = 14'b0000000_0000000;
		Dplus[1495] = 14'b0000000_0000000;
		Dplus[1496] = 14'b0000000_0000000;
		Dplus[1497] = 14'b0000000_0000000;
		Dplus[1498] = 14'b0000000_0000000;
		Dplus[1499] = 14'b0000000_0000000;
		Dplus[1500] = 14'b0000000_0000000;
		Dplus[1501] = 14'b0000000_0000000;
		Dplus[1502] = 14'b0000000_0000000;
		Dplus[1503] = 14'b0000000_0000000;
		Dplus[1504] = 14'b0000000_0000000;
		Dplus[1505] = 14'b0000000_0000000;
		Dplus[1506] = 14'b0000000_0000000;
		Dplus[1507] = 14'b0000000_0000000;
		Dplus[1508] = 14'b0000000_0000000;
		Dplus[1509] = 14'b0000000_0000000;
		Dplus[1510] = 14'b0000000_0000000;
		Dplus[1511] = 14'b0000000_0000000;
		Dplus[1512] = 14'b0000000_0000000;
		Dplus[1513] = 14'b0000000_0000000;
		Dplus[1514] = 14'b0000000_0000000;
		Dplus[1515] = 14'b0000000_0000000;
		Dplus[1516] = 14'b0000000_0000000;
		Dplus[1517] = 14'b0000000_0000000;
		Dplus[1518] = 14'b0000000_0000000;
		Dplus[1519] = 14'b0000000_0000000;
		Dplus[1520] = 14'b0000000_0000000;
		Dplus[1521] = 14'b0000000_0000000;
		Dplus[1522] = 14'b0000000_0000000;
		Dplus[1523] = 14'b0000000_0000000;
		Dplus[1524] = 14'b0000000_0000000;
		Dplus[1525] = 14'b0000000_0000000;
		Dplus[1526] = 14'b0000000_0000000;
		Dplus[1527] = 14'b0000000_0000000;
		Dplus[1528] = 14'b0000000_0000000;
		Dplus[1529] = 14'b0000000_0000000;
		Dplus[1530] = 14'b0000000_0000000;
		Dplus[1531] = 14'b0000000_0000000;
		Dplus[1532] = 14'b0000000_0000000;
		Dplus[1533] = 14'b0000000_0000000;
		Dplus[1534] = 14'b0000000_0000000;
		Dplus[1535] = 14'b0000000_0000000;
		Dplus[1536] = 14'b0000000_0000000;
		Dplus[1537] = 14'b0000000_0000000;
		Dplus[1538] = 14'b0000000_0000000;
		Dplus[1539] = 14'b0000000_0000000;
		Dplus[1540] = 14'b0000000_0000000;
		Dplus[1541] = 14'b0000000_0000000;
		Dplus[1542] = 14'b0000000_0000000;
		Dplus[1543] = 14'b0000000_0000000;
		Dplus[1544] = 14'b0000000_0000000;
		Dplus[1545] = 14'b0000000_0000000;
		Dplus[1546] = 14'b0000000_0000000;
		Dplus[1547] = 14'b0000000_0000000;
		Dplus[1548] = 14'b0000000_0000000;
		Dplus[1549] = 14'b0000000_0000000;
		Dplus[1550] = 14'b0000000_0000000;
		Dplus[1551] = 14'b0000000_0000000;
		Dplus[1552] = 14'b0000000_0000000;
		Dplus[1553] = 14'b0000000_0000000;
		Dplus[1554] = 14'b0000000_0000000;
		Dplus[1555] = 14'b0000000_0000000;
		Dplus[1556] = 14'b0000000_0000000;
		Dplus[1557] = 14'b0000000_0000000;
		Dplus[1558] = 14'b0000000_0000000;
		Dplus[1559] = 14'b0000000_0000000;
		Dplus[1560] = 14'b0000000_0000000;
		Dplus[1561] = 14'b0000000_0000000;
		Dplus[1562] = 14'b0000000_0000000;
		Dplus[1563] = 14'b0000000_0000000;
		Dplus[1564] = 14'b0000000_0000000;
		Dplus[1565] = 14'b0000000_0000000;
		Dplus[1566] = 14'b0000000_0000000;
		Dplus[1567] = 14'b0000000_0000000;
		Dplus[1568] = 14'b0000000_0000000;
		Dplus[1569] = 14'b0000000_0000000;
		Dplus[1570] = 14'b0000000_0000000;
		Dplus[1571] = 14'b0000000_0000000;
		Dplus[1572] = 14'b0000000_0000000;
		Dplus[1573] = 14'b0000000_0000000;
		Dplus[1574] = 14'b0000000_0000000;
		Dplus[1575] = 14'b0000000_0000000;
		Dplus[1576] = 14'b0000000_0000000;
		Dplus[1577] = 14'b0000000_0000000;
		Dplus[1578] = 14'b0000000_0000000;
		Dplus[1579] = 14'b0000000_0000000;
		Dplus[1580] = 14'b0000000_0000000;
		Dplus[1581] = 14'b0000000_0000000;
		Dplus[1582] = 14'b0000000_0000000;
		Dplus[1583] = 14'b0000000_0000000;
		Dplus[1584] = 14'b0000000_0000000;
		Dplus[1585] = 14'b0000000_0000000;
		Dplus[1586] = 14'b0000000_0000000;
		Dplus[1587] = 14'b0000000_0000000;
		Dplus[1588] = 14'b0000000_0000000;
		Dplus[1589] = 14'b0000000_0000000;
		Dplus[1590] = 14'b0000000_0000000;
		Dplus[1591] = 14'b0000000_0000000;
		Dplus[1592] = 14'b0000000_0000000;
		Dplus[1593] = 14'b0000000_0000000;
		Dplus[1594] = 14'b0000000_0000000;
		Dplus[1595] = 14'b0000000_0000000;
		Dplus[1596] = 14'b0000000_0000000;
		Dplus[1597] = 14'b0000000_0000000;
		Dplus[1598] = 14'b0000000_0000000;
		Dplus[1599] = 14'b0000000_0000000;
		Dplus[1600] = 14'b0000000_0000000;
		Dplus[1601] = 14'b0000000_0000000;
		Dplus[1602] = 14'b0000000_0000000;
		Dplus[1603] = 14'b0000000_0000000;
		Dplus[1604] = 14'b0000000_0000000;
		Dplus[1605] = 14'b0000000_0000000;
		Dplus[1606] = 14'b0000000_0000000;
		Dplus[1607] = 14'b0000000_0000000;
		Dplus[1608] = 14'b0000000_0000000;
		Dplus[1609] = 14'b0000000_0000000;
		Dplus[1610] = 14'b0000000_0000000;
		Dplus[1611] = 14'b0000000_0000000;
		Dplus[1612] = 14'b0000000_0000000;
		Dplus[1613] = 14'b0000000_0000000;
		Dplus[1614] = 14'b0000000_0000000;
		Dplus[1615] = 14'b0000000_0000000;
		Dplus[1616] = 14'b0000000_0000000;
		Dplus[1617] = 14'b0000000_0000000;
		Dplus[1618] = 14'b0000000_0000000;
		Dplus[1619] = 14'b0000000_0000000;
		Dplus[1620] = 14'b0000000_0000000;
		Dplus[1621] = 14'b0000000_0000000;
		Dplus[1622] = 14'b0000000_0000000;
		Dplus[1623] = 14'b0000000_0000000;
		Dplus[1624] = 14'b0000000_0000000;
		Dplus[1625] = 14'b0000000_0000000;
		Dplus[1626] = 14'b0000000_0000000;
		Dplus[1627] = 14'b0000000_0000000;
		Dplus[1628] = 14'b0000000_0000000;
		Dplus[1629] = 14'b0000000_0000000;
		Dplus[1630] = 14'b0000000_0000000;
		Dplus[1631] = 14'b0000000_0000000;
		Dplus[1632] = 14'b0000000_0000000;
		Dplus[1633] = 14'b0000000_0000000;
		Dplus[1634] = 14'b0000000_0000000;
		Dplus[1635] = 14'b0000000_0000000;
		Dplus[1636] = 14'b0000000_0000000;
		Dplus[1637] = 14'b0000000_0000000;
		Dplus[1638] = 14'b0000000_0000000;
		Dplus[1639] = 14'b0000000_0000000;
		Dplus[1640] = 14'b0000000_0000000;
		Dplus[1641] = 14'b0000000_0000000;
		Dplus[1642] = 14'b0000000_0000000;
		Dplus[1643] = 14'b0000000_0000000;
		Dplus[1644] = 14'b0000000_0000000;
		Dplus[1645] = 14'b0000000_0000000;
		Dplus[1646] = 14'b0000000_0000000;
		Dplus[1647] = 14'b0000000_0000000;
		Dplus[1648] = 14'b0000000_0000000;
		Dplus[1649] = 14'b0000000_0000000;
		Dplus[1650] = 14'b0000000_0000000;
		Dplus[1651] = 14'b0000000_0000000;
		Dplus[1652] = 14'b0000000_0000000;
		Dplus[1653] = 14'b0000000_0000000;
		Dplus[1654] = 14'b0000000_0000000;
		Dplus[1655] = 14'b0000000_0000000;
		Dplus[1656] = 14'b0000000_0000000;
		Dplus[1657] = 14'b0000000_0000000;
		Dplus[1658] = 14'b0000000_0000000;
		Dplus[1659] = 14'b0000000_0000000;
		Dplus[1660] = 14'b0000000_0000000;
		Dplus[1661] = 14'b0000000_0000000;
		Dplus[1662] = 14'b0000000_0000000;
		Dplus[1663] = 14'b0000000_0000000;
		Dplus[1664] = 14'b0000000_0000000;
		Dplus[1665] = 14'b0000000_0000000;
		Dplus[1666] = 14'b0000000_0000000;
		Dplus[1667] = 14'b0000000_0000000;
		Dplus[1668] = 14'b0000000_0000000;
		Dplus[1669] = 14'b0000000_0000000;
		Dplus[1670] = 14'b0000000_0000000;
		Dplus[1671] = 14'b0000000_0000000;
		Dplus[1672] = 14'b0000000_0000000;
		Dplus[1673] = 14'b0000000_0000000;
		Dplus[1674] = 14'b0000000_0000000;
		Dplus[1675] = 14'b0000000_0000000;
		Dplus[1676] = 14'b0000000_0000000;
		Dplus[1677] = 14'b0000000_0000000;
		Dplus[1678] = 14'b0000000_0000000;
		Dplus[1679] = 14'b0000000_0000000;
		Dplus[1680] = 14'b0000000_0000000;
		Dplus[1681] = 14'b0000000_0000000;
		Dplus[1682] = 14'b0000000_0000000;
		Dplus[1683] = 14'b0000000_0000000;
		Dplus[1684] = 14'b0000000_0000000;
		Dplus[1685] = 14'b0000000_0000000;
		Dplus[1686] = 14'b0000000_0000000;
		Dplus[1687] = 14'b0000000_0000000;
		Dplus[1688] = 14'b0000000_0000000;
		Dplus[1689] = 14'b0000000_0000000;
		Dplus[1690] = 14'b0000000_0000000;
		Dplus[1691] = 14'b0000000_0000000;
		Dplus[1692] = 14'b0000000_0000000;
		Dplus[1693] = 14'b0000000_0000000;
		Dplus[1694] = 14'b0000000_0000000;
		Dplus[1695] = 14'b0000000_0000000;
		Dplus[1696] = 14'b0000000_0000000;
		Dplus[1697] = 14'b0000000_0000000;
		Dplus[1698] = 14'b0000000_0000000;
		Dplus[1699] = 14'b0000000_0000000;
		Dplus[1700] = 14'b0000000_0000000;
		Dplus[1701] = 14'b0000000_0000000;
		Dplus[1702] = 14'b0000000_0000000;
		Dplus[1703] = 14'b0000000_0000000;
		Dplus[1704] = 14'b0000000_0000000;
		Dplus[1705] = 14'b0000000_0000000;
		Dplus[1706] = 14'b0000000_0000000;
		Dplus[1707] = 14'b0000000_0000000;
		Dplus[1708] = 14'b0000000_0000000;
		Dplus[1709] = 14'b0000000_0000000;
		Dplus[1710] = 14'b0000000_0000000;
		Dplus[1711] = 14'b0000000_0000000;
		Dplus[1712] = 14'b0000000_0000000;
		Dplus[1713] = 14'b0000000_0000000;
		Dplus[1714] = 14'b0000000_0000000;
		Dplus[1715] = 14'b0000000_0000000;
		Dplus[1716] = 14'b0000000_0000000;
		Dplus[1717] = 14'b0000000_0000000;
		Dplus[1718] = 14'b0000000_0000000;
		Dplus[1719] = 14'b0000000_0000000;
		Dplus[1720] = 14'b0000000_0000000;
		Dplus[1721] = 14'b0000000_0000000;
		Dplus[1722] = 14'b0000000_0000000;
		Dplus[1723] = 14'b0000000_0000000;
		Dplus[1724] = 14'b0000000_0000000;
		Dplus[1725] = 14'b0000000_0000000;
		Dplus[1726] = 14'b0000000_0000000;
		Dplus[1727] = 14'b0000000_0000000;
		Dplus[1728] = 14'b0000000_0000000;
		Dplus[1729] = 14'b0000000_0000000;
		Dplus[1730] = 14'b0000000_0000000;
		Dplus[1731] = 14'b0000000_0000000;
		Dplus[1732] = 14'b0000000_0000000;
		Dplus[1733] = 14'b0000000_0000000;
		Dplus[1734] = 14'b0000000_0000000;
		Dplus[1735] = 14'b0000000_0000000;
		Dplus[1736] = 14'b0000000_0000000;
		Dplus[1737] = 14'b0000000_0000000;
		Dplus[1738] = 14'b0000000_0000000;
		Dplus[1739] = 14'b0000000_0000000;
		Dplus[1740] = 14'b0000000_0000000;
		Dplus[1741] = 14'b0000000_0000000;
		Dplus[1742] = 14'b0000000_0000000;
		Dplus[1743] = 14'b0000000_0000000;
		Dplus[1744] = 14'b0000000_0000000;
		Dplus[1745] = 14'b0000000_0000000;
		Dplus[1746] = 14'b0000000_0000000;
		Dplus[1747] = 14'b0000000_0000000;
		Dplus[1748] = 14'b0000000_0000000;
		Dplus[1749] = 14'b0000000_0000000;
		Dplus[1750] = 14'b0000000_0000000;
		Dplus[1751] = 14'b0000000_0000000;
		Dplus[1752] = 14'b0000000_0000000;
		Dplus[1753] = 14'b0000000_0000000;
		Dplus[1754] = 14'b0000000_0000000;
		Dplus[1755] = 14'b0000000_0000000;
		Dplus[1756] = 14'b0000000_0000000;
		Dplus[1757] = 14'b0000000_0000000;
		Dplus[1758] = 14'b0000000_0000000;
		Dplus[1759] = 14'b0000000_0000000;
		Dplus[1760] = 14'b0000000_0000000;
		Dplus[1761] = 14'b0000000_0000000;
		Dplus[1762] = 14'b0000000_0000000;
		Dplus[1763] = 14'b0000000_0000000;
		Dplus[1764] = 14'b0000000_0000000;
		Dplus[1765] = 14'b0000000_0000000;
		Dplus[1766] = 14'b0000000_0000000;
		Dplus[1767] = 14'b0000000_0000000;
		Dplus[1768] = 14'b0000000_0000000;
		Dplus[1769] = 14'b0000000_0000000;
		Dplus[1770] = 14'b0000000_0000000;
		Dplus[1771] = 14'b0000000_0000000;
		Dplus[1772] = 14'b0000000_0000000;
		Dplus[1773] = 14'b0000000_0000000;
		Dplus[1774] = 14'b0000000_0000000;
		Dplus[1775] = 14'b0000000_0000000;
		Dplus[1776] = 14'b0000000_0000000;
		Dplus[1777] = 14'b0000000_0000000;
		Dplus[1778] = 14'b0000000_0000000;
		Dplus[1779] = 14'b0000000_0000000;
		Dplus[1780] = 14'b0000000_0000000;
		Dplus[1781] = 14'b0000000_0000000;
		Dplus[1782] = 14'b0000000_0000000;
		Dplus[1783] = 14'b0000000_0000000;
		Dplus[1784] = 14'b0000000_0000000;
		Dplus[1785] = 14'b0000000_0000000;
		Dplus[1786] = 14'b0000000_0000000;
		Dplus[1787] = 14'b0000000_0000000;
		Dplus[1788] = 14'b0000000_0000000;
		Dplus[1789] = 14'b0000000_0000000;
		Dplus[1790] = 14'b0000000_0000000;
		Dplus[1791] = 14'b0000000_0000000;
		Dplus[1792] = 14'b0000000_0000000;
		Dplus[1793] = 14'b0000000_0000000;
		Dplus[1794] = 14'b0000000_0000000;
		Dplus[1795] = 14'b0000000_0000000;
		Dplus[1796] = 14'b0000000_0000000;
		Dplus[1797] = 14'b0000000_0000000;
		Dplus[1798] = 14'b0000000_0000000;
		Dplus[1799] = 14'b0000000_0000000;
		Dplus[1800] = 14'b0000000_0000000;
		Dplus[1801] = 14'b0000000_0000000;
		Dplus[1802] = 14'b0000000_0000000;
		Dplus[1803] = 14'b0000000_0000000;
		Dplus[1804] = 14'b0000000_0000000;
		Dplus[1805] = 14'b0000000_0000000;
		Dplus[1806] = 14'b0000000_0000000;
		Dplus[1807] = 14'b0000000_0000000;
		Dplus[1808] = 14'b0000000_0000000;
		Dplus[1809] = 14'b0000000_0000000;
		Dplus[1810] = 14'b0000000_0000000;
		Dplus[1811] = 14'b0000000_0000000;
		Dplus[1812] = 14'b0000000_0000000;
		Dplus[1813] = 14'b0000000_0000000;
		Dplus[1814] = 14'b0000000_0000000;
		Dplus[1815] = 14'b0000000_0000000;
		Dplus[1816] = 14'b0000000_0000000;
		Dplus[1817] = 14'b0000000_0000000;
		Dplus[1818] = 14'b0000000_0000000;
		Dplus[1819] = 14'b0000000_0000000;
		Dplus[1820] = 14'b0000000_0000000;
		Dplus[1821] = 14'b0000000_0000000;
		Dplus[1822] = 14'b0000000_0000000;
		Dplus[1823] = 14'b0000000_0000000;
		Dplus[1824] = 14'b0000000_0000000;
		Dplus[1825] = 14'b0000000_0000000;
		Dplus[1826] = 14'b0000000_0000000;
		Dplus[1827] = 14'b0000000_0000000;
		Dplus[1828] = 14'b0000000_0000000;
		Dplus[1829] = 14'b0000000_0000000;
		Dplus[1830] = 14'b0000000_0000000;
		Dplus[1831] = 14'b0000000_0000000;
		Dplus[1832] = 14'b0000000_0000000;
		Dplus[1833] = 14'b0000000_0000000;
		Dplus[1834] = 14'b0000000_0000000;
		Dplus[1835] = 14'b0000000_0000000;
		Dplus[1836] = 14'b0000000_0000000;
		Dplus[1837] = 14'b0000000_0000000;
		Dplus[1838] = 14'b0000000_0000000;
		Dplus[1839] = 14'b0000000_0000000;
		Dplus[1840] = 14'b0000000_0000000;
		Dplus[1841] = 14'b0000000_0000000;
		Dplus[1842] = 14'b0000000_0000000;
		Dplus[1843] = 14'b0000000_0000000;
		Dplus[1844] = 14'b0000000_0000000;
		Dplus[1845] = 14'b0000000_0000000;
		Dplus[1846] = 14'b0000000_0000000;
		Dplus[1847] = 14'b0000000_0000000;
		Dplus[1848] = 14'b0000000_0000000;
		Dplus[1849] = 14'b0000000_0000000;
		Dplus[1850] = 14'b0000000_0000000;
		Dplus[1851] = 14'b0000000_0000000;
		Dplus[1852] = 14'b0000000_0000000;
		Dplus[1853] = 14'b0000000_0000000;
		Dplus[1854] = 14'b0000000_0000000;
		Dplus[1855] = 14'b0000000_0000000;
		Dplus[1856] = 14'b0000000_0000000;
		Dplus[1857] = 14'b0000000_0000000;
		Dplus[1858] = 14'b0000000_0000000;
		Dplus[1859] = 14'b0000000_0000000;
		Dplus[1860] = 14'b0000000_0000000;
		Dplus[1861] = 14'b0000000_0000000;
		Dplus[1862] = 14'b0000000_0000000;
		Dplus[1863] = 14'b0000000_0000000;
		Dplus[1864] = 14'b0000000_0000000;
		Dplus[1865] = 14'b0000000_0000000;
		Dplus[1866] = 14'b0000000_0000000;
		Dplus[1867] = 14'b0000000_0000000;
		Dplus[1868] = 14'b0000000_0000000;
		Dplus[1869] = 14'b0000000_0000000;
		Dplus[1870] = 14'b0000000_0000000;
		Dplus[1871] = 14'b0000000_0000000;
		Dplus[1872] = 14'b0000000_0000000;
		Dplus[1873] = 14'b0000000_0000000;
		Dplus[1874] = 14'b0000000_0000000;
		Dplus[1875] = 14'b0000000_0000000;
		Dplus[1876] = 14'b0000000_0000000;
		Dplus[1877] = 14'b0000000_0000000;
		Dplus[1878] = 14'b0000000_0000000;
		Dplus[1879] = 14'b0000000_0000000;
		Dplus[1880] = 14'b0000000_0000000;
		Dplus[1881] = 14'b0000000_0000000;
		Dplus[1882] = 14'b0000000_0000000;
		Dplus[1883] = 14'b0000000_0000000;
		Dplus[1884] = 14'b0000000_0000000;
		Dplus[1885] = 14'b0000000_0000000;
		Dplus[1886] = 14'b0000000_0000000;
		Dplus[1887] = 14'b0000000_0000000;
		Dplus[1888] = 14'b0000000_0000000;
		Dplus[1889] = 14'b0000000_0000000;
		Dplus[1890] = 14'b0000000_0000000;
		Dplus[1891] = 14'b0000000_0000000;
		Dplus[1892] = 14'b0000000_0000000;
		Dplus[1893] = 14'b0000000_0000000;
		Dplus[1894] = 14'b0000000_0000000;
		Dplus[1895] = 14'b0000000_0000000;
		Dplus[1896] = 14'b0000000_0000000;
		Dplus[1897] = 14'b0000000_0000000;
		Dplus[1898] = 14'b0000000_0000000;
		Dplus[1899] = 14'b0000000_0000000;
		Dplus[1900] = 14'b0000000_0000000;
		Dplus[1901] = 14'b0000000_0000000;
		Dplus[1902] = 14'b0000000_0000000;
		Dplus[1903] = 14'b0000000_0000000;
		Dplus[1904] = 14'b0000000_0000000;
		Dplus[1905] = 14'b0000000_0000000;
		Dplus[1906] = 14'b0000000_0000000;
		Dplus[1907] = 14'b0000000_0000000;
		Dplus[1908] = 14'b0000000_0000000;
		Dplus[1909] = 14'b0000000_0000000;
		Dplus[1910] = 14'b0000000_0000000;
		Dplus[1911] = 14'b0000000_0000000;
		Dplus[1912] = 14'b0000000_0000000;
		Dplus[1913] = 14'b0000000_0000000;
		Dplus[1914] = 14'b0000000_0000000;
		Dplus[1915] = 14'b0000000_0000000;
		Dplus[1916] = 14'b0000000_0000000;
		Dplus[1917] = 14'b0000000_0000000;
		Dplus[1918] = 14'b0000000_0000000;
		Dplus[1919] = 14'b0000000_0000000;
		Dplus[1920] = 14'b0000000_0000000;
		Dplus[1921] = 14'b0000000_0000000;
		Dplus[1922] = 14'b0000000_0000000;
		Dplus[1923] = 14'b0000000_0000000;
		Dplus[1924] = 14'b0000000_0000000;
		Dplus[1925] = 14'b0000000_0000000;
		Dplus[1926] = 14'b0000000_0000000;
		Dplus[1927] = 14'b0000000_0000000;
		Dplus[1928] = 14'b0000000_0000000;
		Dplus[1929] = 14'b0000000_0000000;
		Dplus[1930] = 14'b0000000_0000000;
		Dplus[1931] = 14'b0000000_0000000;
		Dplus[1932] = 14'b0000000_0000000;
		Dplus[1933] = 14'b0000000_0000000;
		Dplus[1934] = 14'b0000000_0000000;
		Dplus[1935] = 14'b0000000_0000000;
		Dplus[1936] = 14'b0000000_0000000;
		Dplus[1937] = 14'b0000000_0000000;
		Dplus[1938] = 14'b0000000_0000000;
		Dplus[1939] = 14'b0000000_0000000;
		Dplus[1940] = 14'b0000000_0000000;
		Dplus[1941] = 14'b0000000_0000000;
		Dplus[1942] = 14'b0000000_0000000;
		Dplus[1943] = 14'b0000000_0000000;
		Dplus[1944] = 14'b0000000_0000000;
		Dplus[1945] = 14'b0000000_0000000;
		Dplus[1946] = 14'b0000000_0000000;
		Dplus[1947] = 14'b0000000_0000000;
		Dplus[1948] = 14'b0000000_0000000;
		Dplus[1949] = 14'b0000000_0000000;
		Dplus[1950] = 14'b0000000_0000000;
		Dplus[1951] = 14'b0000000_0000000;
		Dplus[1952] = 14'b0000000_0000000;
		Dplus[1953] = 14'b0000000_0000000;
		Dplus[1954] = 14'b0000000_0000000;
		Dplus[1955] = 14'b0000000_0000000;
		Dplus[1956] = 14'b0000000_0000000;
		Dplus[1957] = 14'b0000000_0000000;
		Dplus[1958] = 14'b0000000_0000000;
		Dplus[1959] = 14'b0000000_0000000;
		Dplus[1960] = 14'b0000000_0000000;
		Dplus[1961] = 14'b0000000_0000000;
		Dplus[1962] = 14'b0000000_0000000;
		Dplus[1963] = 14'b0000000_0000000;
		Dplus[1964] = 14'b0000000_0000000;
		Dplus[1965] = 14'b0000000_0000000;
		Dplus[1966] = 14'b0000000_0000000;
		Dplus[1967] = 14'b0000000_0000000;
		Dplus[1968] = 14'b0000000_0000000;
		Dplus[1969] = 14'b0000000_0000000;
		Dplus[1970] = 14'b0000000_0000000;
		Dplus[1971] = 14'b0000000_0000000;
		Dplus[1972] = 14'b0000000_0000000;
		Dplus[1973] = 14'b0000000_0000000;
		Dplus[1974] = 14'b0000000_0000000;
		Dplus[1975] = 14'b0000000_0000000;
		Dplus[1976] = 14'b0000000_0000000;
		Dplus[1977] = 14'b0000000_0000000;
		Dplus[1978] = 14'b0000000_0000000;
		Dplus[1979] = 14'b0000000_0000000;
		Dplus[1980] = 14'b0000000_0000000;
		Dplus[1981] = 14'b0000000_0000000;
		Dplus[1982] = 14'b0000000_0000000;
		Dplus[1983] = 14'b0000000_0000000;
		Dplus[1984] = 14'b0000000_0000000;
		Dplus[1985] = 14'b0000000_0000000;
		Dplus[1986] = 14'b0000000_0000000;
		Dplus[1987] = 14'b0000000_0000000;
		Dplus[1988] = 14'b0000000_0000000;
		Dplus[1989] = 14'b0000000_0000000;
		Dplus[1990] = 14'b0000000_0000000;
		Dplus[1991] = 14'b0000000_0000000;
		Dplus[1992] = 14'b0000000_0000000;
		Dplus[1993] = 14'b0000000_0000000;
		Dplus[1994] = 14'b0000000_0000000;
		Dplus[1995] = 14'b0000000_0000000;
		Dplus[1996] = 14'b0000000_0000000;
		Dplus[1997] = 14'b0000000_0000000;
		Dplus[1998] = 14'b0000000_0000000;
		Dplus[1999] = 14'b0000000_0000000;
		Dplus[2000] = 14'b0000000_0000000;
		Dplus[2001] = 14'b0000000_0000000;
		Dplus[2002] = 14'b0000000_0000000;
		Dplus[2003] = 14'b0000000_0000000;
		Dplus[2004] = 14'b0000000_0000000;
		Dplus[2005] = 14'b0000000_0000000;
		Dplus[2006] = 14'b0000000_0000000;
		Dplus[2007] = 14'b0000000_0000000;
		Dplus[2008] = 14'b0000000_0000000;
		Dplus[2009] = 14'b0000000_0000000;
		Dplus[2010] = 14'b0000000_0000000;
		Dplus[2011] = 14'b0000000_0000000;
		Dplus[2012] = 14'b0000000_0000000;
		Dplus[2013] = 14'b0000000_0000000;
		Dplus[2014] = 14'b0000000_0000000;
		Dplus[2015] = 14'b0000000_0000000;
		Dplus[2016] = 14'b0000000_0000000;
		Dplus[2017] = 14'b0000000_0000000;
		Dplus[2018] = 14'b0000000_0000000;
		Dplus[2019] = 14'b0000000_0000000;
		Dplus[2020] = 14'b0000000_0000000;
		Dplus[2021] = 14'b0000000_0000000;
		Dplus[2022] = 14'b0000000_0000000;
		Dplus[2023] = 14'b0000000_0000000;
		Dplus[2024] = 14'b0000000_0000000;
		Dplus[2025] = 14'b0000000_0000000;
		Dplus[2026] = 14'b0000000_0000000;
		Dplus[2027] = 14'b0000000_0000000;
		Dplus[2028] = 14'b0000000_0000000;
		Dplus[2029] = 14'b0000000_0000000;
		Dplus[2030] = 14'b0000000_0000000;
		Dplus[2031] = 14'b0000000_0000000;
		Dplus[2032] = 14'b0000000_0000000;
		Dplus[2033] = 14'b0000000_0000000;
		Dplus[2034] = 14'b0000000_0000000;
		Dplus[2035] = 14'b0000000_0000000;
		Dplus[2036] = 14'b0000000_0000000;
		Dplus[2037] = 14'b0000000_0000000;
		Dplus[2038] = 14'b0000000_0000000;
		Dplus[2039] = 14'b0000000_0000000;
		Dplus[2040] = 14'b0000000_0000000;
		Dplus[2041] = 14'b0000000_0000000;
		Dplus[2042] = 14'b0000000_0000000;
		Dplus[2043] = 14'b0000000_0000000;
		Dplus[2044] = 14'b0000000_0000000;
		Dplus[2045] = 14'b0000000_0000000;
		Dplus[2046] = 14'b0000000_0000000;
		Dplus[2047] = 14'b0000000_0000000;
		Dplus[2048] = 14'b0000000_0000000;
		Dplus[2049] = 14'b0000000_0000000;
		Dplus[2050] = 14'b0000000_0000000;
		Dplus[2051] = 14'b0000000_0000000;
		Dplus[2052] = 14'b0000000_0000000;
		Dplus[2053] = 14'b0000000_0000000;
		Dplus[2054] = 14'b0000000_0000000;
		Dplus[2055] = 14'b0000000_0000000;
		Dplus[2056] = 14'b0000000_0000000;
		Dplus[2057] = 14'b0000000_0000000;
		Dplus[2058] = 14'b0000000_0000000;
		Dplus[2059] = 14'b0000000_0000000;
		Dplus[2060] = 14'b0000000_0000000;
		Dplus[2061] = 14'b0000000_0000000;
		Dplus[2062] = 14'b0000000_0000000;
		Dplus[2063] = 14'b0000000_0000000;
		Dplus[2064] = 14'b0000000_0000000;
		Dplus[2065] = 14'b0000000_0000000;
		Dplus[2066] = 14'b0000000_0000000;
		Dplus[2067] = 14'b0000000_0000000;
		Dplus[2068] = 14'b0000000_0000000;
		Dplus[2069] = 14'b0000000_0000000;
		Dplus[2070] = 14'b0000000_0000000;
		Dplus[2071] = 14'b0000000_0000000;
		Dplus[2072] = 14'b0000000_0000000;
		Dplus[2073] = 14'b0000000_0000000;
		Dplus[2074] = 14'b0000000_0000000;
		Dplus[2075] = 14'b0000000_0000000;
		Dplus[2076] = 14'b0000000_0000000;
		Dplus[2077] = 14'b0000000_0000000;
		Dplus[2078] = 14'b0000000_0000000;
		Dplus[2079] = 14'b0000000_0000000;
		Dplus[2080] = 14'b0000000_0000000;
		Dplus[2081] = 14'b0000000_0000000;
		Dplus[2082] = 14'b0000000_0000000;
		Dplus[2083] = 14'b0000000_0000000;
		Dplus[2084] = 14'b0000000_0000000;
		Dplus[2085] = 14'b0000000_0000000;
		Dplus[2086] = 14'b0000000_0000000;
		Dplus[2087] = 14'b0000000_0000000;
		Dplus[2088] = 14'b0000000_0000000;
		Dplus[2089] = 14'b0000000_0000000;
		Dplus[2090] = 14'b0000000_0000000;
		Dplus[2091] = 14'b0000000_0000000;
		Dplus[2092] = 14'b0000000_0000000;
		Dplus[2093] = 14'b0000000_0000000;
		Dplus[2094] = 14'b0000000_0000000;
		Dplus[2095] = 14'b0000000_0000000;
		Dplus[2096] = 14'b0000000_0000000;
		Dplus[2097] = 14'b0000000_0000000;
		Dplus[2098] = 14'b0000000_0000000;
		Dplus[2099] = 14'b0000000_0000000;
		Dplus[2100] = 14'b0000000_0000000;
		Dplus[2101] = 14'b0000000_0000000;
		Dplus[2102] = 14'b0000000_0000000;
		Dplus[2103] = 14'b0000000_0000000;
		Dplus[2104] = 14'b0000000_0000000;
		Dplus[2105] = 14'b0000000_0000000;
		Dplus[2106] = 14'b0000000_0000000;
		Dplus[2107] = 14'b0000000_0000000;
		Dplus[2108] = 14'b0000000_0000000;
		Dplus[2109] = 14'b0000000_0000000;
		Dplus[2110] = 14'b0000000_0000000;
		Dplus[2111] = 14'b0000000_0000000;
		Dplus[2112] = 14'b0000000_0000000;
		Dplus[2113] = 14'b0000000_0000000;
		Dplus[2114] = 14'b0000000_0000000;
		Dplus[2115] = 14'b0000000_0000000;
		Dplus[2116] = 14'b0000000_0000000;
		Dplus[2117] = 14'b0000000_0000000;
		Dplus[2118] = 14'b0000000_0000000;
		Dplus[2119] = 14'b0000000_0000000;
		Dplus[2120] = 14'b0000000_0000000;
		Dplus[2121] = 14'b0000000_0000000;
		Dplus[2122] = 14'b0000000_0000000;
		Dplus[2123] = 14'b0000000_0000000;
		Dplus[2124] = 14'b0000000_0000000;
		Dplus[2125] = 14'b0000000_0000000;
		Dplus[2126] = 14'b0000000_0000000;
		Dplus[2127] = 14'b0000000_0000000;
		Dplus[2128] = 14'b0000000_0000000;
		Dplus[2129] = 14'b0000000_0000000;
		Dplus[2130] = 14'b0000000_0000000;
		Dplus[2131] = 14'b0000000_0000000;
		Dplus[2132] = 14'b0000000_0000000;
		Dplus[2133] = 14'b0000000_0000000;
		Dplus[2134] = 14'b0000000_0000000;
		Dplus[2135] = 14'b0000000_0000000;
		Dplus[2136] = 14'b0000000_0000000;
		Dplus[2137] = 14'b0000000_0000000;
		Dplus[2138] = 14'b0000000_0000000;
		Dplus[2139] = 14'b0000000_0000000;
		Dplus[2140] = 14'b0000000_0000000;
		Dplus[2141] = 14'b0000000_0000000;
		Dplus[2142] = 14'b0000000_0000000;
		Dplus[2143] = 14'b0000000_0000000;
		Dplus[2144] = 14'b0000000_0000000;
		Dplus[2145] = 14'b0000000_0000000;
		Dplus[2146] = 14'b0000000_0000000;
		Dplus[2147] = 14'b0000000_0000000;
		Dplus[2148] = 14'b0000000_0000000;
		Dplus[2149] = 14'b0000000_0000000;
		Dplus[2150] = 14'b0000000_0000000;
		Dplus[2151] = 14'b0000000_0000000;
		Dplus[2152] = 14'b0000000_0000000;
		Dplus[2153] = 14'b0000000_0000000;
		Dplus[2154] = 14'b0000000_0000000;
		Dplus[2155] = 14'b0000000_0000000;
		Dplus[2156] = 14'b0000000_0000000;
		Dplus[2157] = 14'b0000000_0000000;
		Dplus[2158] = 14'b0000000_0000000;
		Dplus[2159] = 14'b0000000_0000000;
		Dplus[2160] = 14'b0000000_0000000;
		Dplus[2161] = 14'b0000000_0000000;
		Dplus[2162] = 14'b0000000_0000000;
		Dplus[2163] = 14'b0000000_0000000;
		Dplus[2164] = 14'b0000000_0000000;
		Dplus[2165] = 14'b0000000_0000000;
		Dplus[2166] = 14'b0000000_0000000;
		Dplus[2167] = 14'b0000000_0000000;
		Dplus[2168] = 14'b0000000_0000000;
		Dplus[2169] = 14'b0000000_0000000;
		Dplus[2170] = 14'b0000000_0000000;
		Dplus[2171] = 14'b0000000_0000000;
		Dplus[2172] = 14'b0000000_0000000;
		Dplus[2173] = 14'b0000000_0000000;
		Dplus[2174] = 14'b0000000_0000000;
		Dplus[2175] = 14'b0000000_0000000;
		Dplus[2176] = 14'b0000000_0000000;
		Dplus[2177] = 14'b0000000_0000000;
		Dplus[2178] = 14'b0000000_0000000;
		Dplus[2179] = 14'b0000000_0000000;
		Dplus[2180] = 14'b0000000_0000000;
		Dplus[2181] = 14'b0000000_0000000;
		Dplus[2182] = 14'b0000000_0000000;
		Dplus[2183] = 14'b0000000_0000000;
		Dplus[2184] = 14'b0000000_0000000;
		Dplus[2185] = 14'b0000000_0000000;
		Dplus[2186] = 14'b0000000_0000000;
		Dplus[2187] = 14'b0000000_0000000;
		Dplus[2188] = 14'b0000000_0000000;
		Dplus[2189] = 14'b0000000_0000000;
		Dplus[2190] = 14'b0000000_0000000;
		Dplus[2191] = 14'b0000000_0000000;
		Dplus[2192] = 14'b0000000_0000000;
		Dplus[2193] = 14'b0000000_0000000;
		Dplus[2194] = 14'b0000000_0000000;
		Dplus[2195] = 14'b0000000_0000000;
		Dplus[2196] = 14'b0000000_0000000;
		Dplus[2197] = 14'b0000000_0000000;
		Dplus[2198] = 14'b0000000_0000000;
		Dplus[2199] = 14'b0000000_0000000;
		Dplus[2200] = 14'b0000000_0000000;
		Dplus[2201] = 14'b0000000_0000000;
		Dplus[2202] = 14'b0000000_0000000;
		Dplus[2203] = 14'b0000000_0000000;
		Dplus[2204] = 14'b0000000_0000000;
		Dplus[2205] = 14'b0000000_0000000;
		Dplus[2206] = 14'b0000000_0000000;
		Dplus[2207] = 14'b0000000_0000000;
		Dplus[2208] = 14'b0000000_0000000;
		Dplus[2209] = 14'b0000000_0000000;
		Dplus[2210] = 14'b0000000_0000000;
		Dplus[2211] = 14'b0000000_0000000;
		Dplus[2212] = 14'b0000000_0000000;
		Dplus[2213] = 14'b0000000_0000000;
		Dplus[2214] = 14'b0000000_0000000;
		Dplus[2215] = 14'b0000000_0000000;
		Dplus[2216] = 14'b0000000_0000000;
		Dplus[2217] = 14'b0000000_0000000;
		Dplus[2218] = 14'b0000000_0000000;
		Dplus[2219] = 14'b0000000_0000000;
		Dplus[2220] = 14'b0000000_0000000;
		Dplus[2221] = 14'b0000000_0000000;
		Dplus[2222] = 14'b0000000_0000000;
		Dplus[2223] = 14'b0000000_0000000;
		Dplus[2224] = 14'b0000000_0000000;
		Dplus[2225] = 14'b0000000_0000000;
		Dplus[2226] = 14'b0000000_0000000;
		Dplus[2227] = 14'b0000000_0000000;
		Dplus[2228] = 14'b0000000_0000000;
		Dplus[2229] = 14'b0000000_0000000;
		Dplus[2230] = 14'b0000000_0000000;
		Dplus[2231] = 14'b0000000_0000000;
		Dplus[2232] = 14'b0000000_0000000;
		Dplus[2233] = 14'b0000000_0000000;
		Dplus[2234] = 14'b0000000_0000000;
		Dplus[2235] = 14'b0000000_0000000;
		Dplus[2236] = 14'b0000000_0000000;
		Dplus[2237] = 14'b0000000_0000000;
		Dplus[2238] = 14'b0000000_0000000;
		Dplus[2239] = 14'b0000000_0000000;
		Dplus[2240] = 14'b0000000_0000000;
		Dplus[2241] = 14'b0000000_0000000;
		Dplus[2242] = 14'b0000000_0000000;
		Dplus[2243] = 14'b0000000_0000000;
		Dplus[2244] = 14'b0000000_0000000;
		Dplus[2245] = 14'b0000000_0000000;
		Dplus[2246] = 14'b0000000_0000000;
		Dplus[2247] = 14'b0000000_0000000;
		Dplus[2248] = 14'b0000000_0000000;
		Dplus[2249] = 14'b0000000_0000000;
		Dplus[2250] = 14'b0000000_0000000;
		Dplus[2251] = 14'b0000000_0000000;
		Dplus[2252] = 14'b0000000_0000000;
		Dplus[2253] = 14'b0000000_0000000;
		Dplus[2254] = 14'b0000000_0000000;
		Dplus[2255] = 14'b0000000_0000000;
		Dplus[2256] = 14'b0000000_0000000;
		Dplus[2257] = 14'b0000000_0000000;
		Dplus[2258] = 14'b0000000_0000000;
		Dplus[2259] = 14'b0000000_0000000;
		Dplus[2260] = 14'b0000000_0000000;
		Dplus[2261] = 14'b0000000_0000000;
		Dplus[2262] = 14'b0000000_0000000;
		Dplus[2263] = 14'b0000000_0000000;
		Dplus[2264] = 14'b0000000_0000000;
		Dplus[2265] = 14'b0000000_0000000;
		Dplus[2266] = 14'b0000000_0000000;
		Dplus[2267] = 14'b0000000_0000000;
		Dplus[2268] = 14'b0000000_0000000;
		Dplus[2269] = 14'b0000000_0000000;
		Dplus[2270] = 14'b0000000_0000000;
		Dplus[2271] = 14'b0000000_0000000;
		Dplus[2272] = 14'b0000000_0000000;
		Dplus[2273] = 14'b0000000_0000000;
		Dplus[2274] = 14'b0000000_0000000;
		Dplus[2275] = 14'b0000000_0000000;
		Dplus[2276] = 14'b0000000_0000000;
		Dplus[2277] = 14'b0000000_0000000;
		Dplus[2278] = 14'b0000000_0000000;
		Dplus[2279] = 14'b0000000_0000000;
		Dplus[2280] = 14'b0000000_0000000;
		Dplus[2281] = 14'b0000000_0000000;
		Dplus[2282] = 14'b0000000_0000000;
		Dplus[2283] = 14'b0000000_0000000;
		Dplus[2284] = 14'b0000000_0000000;
		Dplus[2285] = 14'b0000000_0000000;
		Dplus[2286] = 14'b0000000_0000000;
		Dplus[2287] = 14'b0000000_0000000;
		Dplus[2288] = 14'b0000000_0000000;
		Dplus[2289] = 14'b0000000_0000000;
		Dplus[2290] = 14'b0000000_0000000;
		Dplus[2291] = 14'b0000000_0000000;
		Dplus[2292] = 14'b0000000_0000000;
		Dplus[2293] = 14'b0000000_0000000;
		Dplus[2294] = 14'b0000000_0000000;
		Dplus[2295] = 14'b0000000_0000000;
		Dplus[2296] = 14'b0000000_0000000;
		Dplus[2297] = 14'b0000000_0000000;
		Dplus[2298] = 14'b0000000_0000000;
		Dplus[2299] = 14'b0000000_0000000;
		Dplus[2300] = 14'b0000000_0000000;
		Dplus[2301] = 14'b0000000_0000000;
		Dplus[2302] = 14'b0000000_0000000;
		Dplus[2303] = 14'b0000000_0000000;
		Dplus[2304] = 14'b0000000_0000000;
		Dplus[2305] = 14'b0000000_0000000;
		Dplus[2306] = 14'b0000000_0000000;
		Dplus[2307] = 14'b0000000_0000000;
		Dplus[2308] = 14'b0000000_0000000;
		Dplus[2309] = 14'b0000000_0000000;
		Dplus[2310] = 14'b0000000_0000000;
		Dplus[2311] = 14'b0000000_0000000;
		Dplus[2312] = 14'b0000000_0000000;
		Dplus[2313] = 14'b0000000_0000000;
		Dplus[2314] = 14'b0000000_0000000;
		Dplus[2315] = 14'b0000000_0000000;
		Dplus[2316] = 14'b0000000_0000000;
		Dplus[2317] = 14'b0000000_0000000;
		Dplus[2318] = 14'b0000000_0000000;
		Dplus[2319] = 14'b0000000_0000000;
		Dplus[2320] = 14'b0000000_0000000;
		Dplus[2321] = 14'b0000000_0000000;
		Dplus[2322] = 14'b0000000_0000000;
		Dplus[2323] = 14'b0000000_0000000;
		Dplus[2324] = 14'b0000000_0000000;
		Dplus[2325] = 14'b0000000_0000000;
		Dplus[2326] = 14'b0000000_0000000;
		Dplus[2327] = 14'b0000000_0000000;
		Dplus[2328] = 14'b0000000_0000000;
		Dplus[2329] = 14'b0000000_0000000;
		Dplus[2330] = 14'b0000000_0000000;
		Dplus[2331] = 14'b0000000_0000000;
		Dplus[2332] = 14'b0000000_0000000;
		Dplus[2333] = 14'b0000000_0000000;
		Dplus[2334] = 14'b0000000_0000000;
		Dplus[2335] = 14'b0000000_0000000;
		Dplus[2336] = 14'b0000000_0000000;
		Dplus[2337] = 14'b0000000_0000000;
		Dplus[2338] = 14'b0000000_0000000;
		Dplus[2339] = 14'b0000000_0000000;
		Dplus[2340] = 14'b0000000_0000000;
		Dplus[2341] = 14'b0000000_0000000;
		Dplus[2342] = 14'b0000000_0000000;
		Dplus[2343] = 14'b0000000_0000000;
		Dplus[2344] = 14'b0000000_0000000;
		Dplus[2345] = 14'b0000000_0000000;
		Dplus[2346] = 14'b0000000_0000000;
		Dplus[2347] = 14'b0000000_0000000;
		Dplus[2348] = 14'b0000000_0000000;
		Dplus[2349] = 14'b0000000_0000000;
		Dplus[2350] = 14'b0000000_0000000;
		Dplus[2351] = 14'b0000000_0000000;
		Dplus[2352] = 14'b0000000_0000000;
		Dplus[2353] = 14'b0000000_0000000;
		Dplus[2354] = 14'b0000000_0000000;
		Dplus[2355] = 14'b0000000_0000000;
		Dplus[2356] = 14'b0000000_0000000;
		Dplus[2357] = 14'b0000000_0000000;
		Dplus[2358] = 14'b0000000_0000000;
		Dplus[2359] = 14'b0000000_0000000;
		Dplus[2360] = 14'b0000000_0000000;
		Dplus[2361] = 14'b0000000_0000000;
		Dplus[2362] = 14'b0000000_0000000;
		Dplus[2363] = 14'b0000000_0000000;
		Dplus[2364] = 14'b0000000_0000000;
		Dplus[2365] = 14'b0000000_0000000;
		Dplus[2366] = 14'b0000000_0000000;
		Dplus[2367] = 14'b0000000_0000000;
		Dplus[2368] = 14'b0000000_0000000;
		Dplus[2369] = 14'b0000000_0000000;
		Dplus[2370] = 14'b0000000_0000000;
		Dplus[2371] = 14'b0000000_0000000;
		Dplus[2372] = 14'b0000000_0000000;
		Dplus[2373] = 14'b0000000_0000000;
		Dplus[2374] = 14'b0000000_0000000;
		Dplus[2375] = 14'b0000000_0000000;
		Dplus[2376] = 14'b0000000_0000000;
		Dplus[2377] = 14'b0000000_0000000;
		Dplus[2378] = 14'b0000000_0000000;
		Dplus[2379] = 14'b0000000_0000000;
		Dplus[2380] = 14'b0000000_0000000;
		Dplus[2381] = 14'b0000000_0000000;
		Dplus[2382] = 14'b0000000_0000000;
		Dplus[2383] = 14'b0000000_0000000;
		Dplus[2384] = 14'b0000000_0000000;
		Dplus[2385] = 14'b0000000_0000000;
		Dplus[2386] = 14'b0000000_0000000;
		Dplus[2387] = 14'b0000000_0000000;
		Dplus[2388] = 14'b0000000_0000000;
		Dplus[2389] = 14'b0000000_0000000;
		Dplus[2390] = 14'b0000000_0000000;
		Dplus[2391] = 14'b0000000_0000000;
		Dplus[2392] = 14'b0000000_0000000;
		Dplus[2393] = 14'b0000000_0000000;
		Dplus[2394] = 14'b0000000_0000000;
		Dplus[2395] = 14'b0000000_0000000;
		Dplus[2396] = 14'b0000000_0000000;
		Dplus[2397] = 14'b0000000_0000000;
		Dplus[2398] = 14'b0000000_0000000;
		Dplus[2399] = 14'b0000000_0000000;
		Dplus[2400] = 14'b0000000_0000000;
		Dplus[2401] = 14'b0000000_0000000;
		Dplus[2402] = 14'b0000000_0000000;
		Dplus[2403] = 14'b0000000_0000000;
		Dplus[2404] = 14'b0000000_0000000;
		Dplus[2405] = 14'b0000000_0000000;
		Dplus[2406] = 14'b0000000_0000000;
		Dplus[2407] = 14'b0000000_0000000;
		Dplus[2408] = 14'b0000000_0000000;
		Dplus[2409] = 14'b0000000_0000000;
		Dplus[2410] = 14'b0000000_0000000;
		Dplus[2411] = 14'b0000000_0000000;
		Dplus[2412] = 14'b0000000_0000000;
		Dplus[2413] = 14'b0000000_0000000;
		Dplus[2414] = 14'b0000000_0000000;
		Dplus[2415] = 14'b0000000_0000000;
		Dplus[2416] = 14'b0000000_0000000;
		Dplus[2417] = 14'b0000000_0000000;
		Dplus[2418] = 14'b0000000_0000000;
		Dplus[2419] = 14'b0000000_0000000;
		Dplus[2420] = 14'b0000000_0000000;
		Dplus[2421] = 14'b0000000_0000000;
		Dplus[2422] = 14'b0000000_0000000;
		Dplus[2423] = 14'b0000000_0000000;
		Dplus[2424] = 14'b0000000_0000000;
		Dplus[2425] = 14'b0000000_0000000;
		Dplus[2426] = 14'b0000000_0000000;
		Dplus[2427] = 14'b0000000_0000000;
		Dplus[2428] = 14'b0000000_0000000;
		Dplus[2429] = 14'b0000000_0000000;
		Dplus[2430] = 14'b0000000_0000000;
		Dplus[2431] = 14'b0000000_0000000;
		Dplus[2432] = 14'b0000000_0000000;
		Dplus[2433] = 14'b0000000_0000000;
		Dplus[2434] = 14'b0000000_0000000;
		Dplus[2435] = 14'b0000000_0000000;
		Dplus[2436] = 14'b0000000_0000000;
		Dplus[2437] = 14'b0000000_0000000;
		Dplus[2438] = 14'b0000000_0000000;
		Dplus[2439] = 14'b0000000_0000000;
		Dplus[2440] = 14'b0000000_0000000;
		Dplus[2441] = 14'b0000000_0000000;
		Dplus[2442] = 14'b0000000_0000000;
		Dplus[2443] = 14'b0000000_0000000;
		Dplus[2444] = 14'b0000000_0000000;
		Dplus[2445] = 14'b0000000_0000000;
		Dplus[2446] = 14'b0000000_0000000;
		Dplus[2447] = 14'b0000000_0000000;
		Dplus[2448] = 14'b0000000_0000000;
		Dplus[2449] = 14'b0000000_0000000;
		Dplus[2450] = 14'b0000000_0000000;
		Dplus[2451] = 14'b0000000_0000000;
		Dplus[2452] = 14'b0000000_0000000;
		Dplus[2453] = 14'b0000000_0000000;
		Dplus[2454] = 14'b0000000_0000000;
		Dplus[2455] = 14'b0000000_0000000;
		Dplus[2456] = 14'b0000000_0000000;
		Dplus[2457] = 14'b0000000_0000000;
		Dplus[2458] = 14'b0000000_0000000;
		Dplus[2459] = 14'b0000000_0000000;
		Dplus[2460] = 14'b0000000_0000000;
		Dplus[2461] = 14'b0000000_0000000;
		Dplus[2462] = 14'b0000000_0000000;
		Dplus[2463] = 14'b0000000_0000000;
		Dplus[2464] = 14'b0000000_0000000;
		Dplus[2465] = 14'b0000000_0000000;
		Dplus[2466] = 14'b0000000_0000000;
		Dplus[2467] = 14'b0000000_0000000;
		Dplus[2468] = 14'b0000000_0000000;
		Dplus[2469] = 14'b0000000_0000000;
		Dplus[2470] = 14'b0000000_0000000;
		Dplus[2471] = 14'b0000000_0000000;
		Dplus[2472] = 14'b0000000_0000000;
		Dplus[2473] = 14'b0000000_0000000;
		Dplus[2474] = 14'b0000000_0000000;
		Dplus[2475] = 14'b0000000_0000000;
		Dplus[2476] = 14'b0000000_0000000;
		Dplus[2477] = 14'b0000000_0000000;
		Dplus[2478] = 14'b0000000_0000000;
		Dplus[2479] = 14'b0000000_0000000;
		Dplus[2480] = 14'b0000000_0000000;
		Dplus[2481] = 14'b0000000_0000000;
		Dplus[2482] = 14'b0000000_0000000;
		Dplus[2483] = 14'b0000000_0000000;
		Dplus[2484] = 14'b0000000_0000000;
		Dplus[2485] = 14'b0000000_0000000;
		Dplus[2486] = 14'b0000000_0000000;
		Dplus[2487] = 14'b0000000_0000000;
		Dplus[2488] = 14'b0000000_0000000;
		Dplus[2489] = 14'b0000000_0000000;
		Dplus[2490] = 14'b0000000_0000000;
		Dplus[2491] = 14'b0000000_0000000;
		Dplus[2492] = 14'b0000000_0000000;
		Dplus[2493] = 14'b0000000_0000000;
		Dplus[2494] = 14'b0000000_0000000;
		Dplus[2495] = 14'b0000000_0000000;
		Dplus[2496] = 14'b0000000_0000000;
		Dplus[2497] = 14'b0000000_0000000;
		Dplus[2498] = 14'b0000000_0000000;
		Dplus[2499] = 14'b0000000_0000000;
		Dplus[2500] = 14'b0000000_0000000;
		Dplus[2501] = 14'b0000000_0000000;
		Dplus[2502] = 14'b0000000_0000000;
		Dplus[2503] = 14'b0000000_0000000;
		Dplus[2504] = 14'b0000000_0000000;
		Dplus[2505] = 14'b0000000_0000000;
		Dplus[2506] = 14'b0000000_0000000;
		Dplus[2507] = 14'b0000000_0000000;
		Dplus[2508] = 14'b0000000_0000000;
		Dplus[2509] = 14'b0000000_0000000;
		Dplus[2510] = 14'b0000000_0000000;
		Dplus[2511] = 14'b0000000_0000000;
		Dplus[2512] = 14'b0000000_0000000;
		Dplus[2513] = 14'b0000000_0000000;
		Dplus[2514] = 14'b0000000_0000000;
		Dplus[2515] = 14'b0000000_0000000;
		Dplus[2516] = 14'b0000000_0000000;
		Dplus[2517] = 14'b0000000_0000000;
		Dplus[2518] = 14'b0000000_0000000;
		Dplus[2519] = 14'b0000000_0000000;
		Dplus[2520] = 14'b0000000_0000000;
		Dplus[2521] = 14'b0000000_0000000;
		Dplus[2522] = 14'b0000000_0000000;
		Dplus[2523] = 14'b0000000_0000000;
		Dplus[2524] = 14'b0000000_0000000;
		Dplus[2525] = 14'b0000000_0000000;
		Dplus[2526] = 14'b0000000_0000000;
		Dplus[2527] = 14'b0000000_0000000;
		Dplus[2528] = 14'b0000000_0000000;
		Dplus[2529] = 14'b0000000_0000000;
		Dplus[2530] = 14'b0000000_0000000;
		Dplus[2531] = 14'b0000000_0000000;
		Dplus[2532] = 14'b0000000_0000000;
		Dplus[2533] = 14'b0000000_0000000;
		Dplus[2534] = 14'b0000000_0000000;
		Dplus[2535] = 14'b0000000_0000000;
		Dplus[2536] = 14'b0000000_0000000;
		Dplus[2537] = 14'b0000000_0000000;
		Dplus[2538] = 14'b0000000_0000000;
		Dplus[2539] = 14'b0000000_0000000;
		Dplus[2540] = 14'b0000000_0000000;
		Dplus[2541] = 14'b0000000_0000000;
		Dplus[2542] = 14'b0000000_0000000;
		Dplus[2543] = 14'b0000000_0000000;
		Dplus[2544] = 14'b0000000_0000000;
		Dplus[2545] = 14'b0000000_0000000;
		Dplus[2546] = 14'b0000000_0000000;
		Dplus[2547] = 14'b0000000_0000000;
		Dplus[2548] = 14'b0000000_0000000;
		Dplus[2549] = 14'b0000000_0000000;
		Dplus[2550] = 14'b0000000_0000000;
		Dplus[2551] = 14'b0000000_0000000;
		Dplus[2552] = 14'b0000000_0000000;
		Dplus[2553] = 14'b0000000_0000000;
		Dplus[2554] = 14'b0000000_0000000;
		Dplus[2555] = 14'b0000000_0000000;
		Dplus[2556] = 14'b0000000_0000000;
		Dplus[2557] = 14'b0000000_0000000;
		Dplus[2558] = 14'b0000000_0000000;
		Dplus[2559] = 14'b0000000_0000000;
		Dplus[2560] = 14'b0000000_0000000;
		Dplus[2561] = 14'b0000000_0000000;
		Dplus[2562] = 14'b0000000_0000000;
		Dplus[2563] = 14'b0000000_0000000;
		Dplus[2564] = 14'b0000000_0000000;
		Dplus[2565] = 14'b0000000_0000000;
		Dplus[2566] = 14'b0000000_0000000;
		Dplus[2567] = 14'b0000000_0000000;
		Dplus[2568] = 14'b0000000_0000000;
		Dplus[2569] = 14'b0000000_0000000;
		Dplus[2570] = 14'b0000000_0000000;
		Dplus[2571] = 14'b0000000_0000000;
		Dplus[2572] = 14'b0000000_0000000;
		Dplus[2573] = 14'b0000000_0000000;
		Dplus[2574] = 14'b0000000_0000000;
		Dplus[2575] = 14'b0000000_0000000;
		Dplus[2576] = 14'b0000000_0000000;
		Dplus[2577] = 14'b0000000_0000000;
		Dplus[2578] = 14'b0000000_0000000;
		Dplus[2579] = 14'b0000000_0000000;
		Dplus[2580] = 14'b0000000_0000000;
		Dplus[2581] = 14'b0000000_0000000;
		Dplus[2582] = 14'b0000000_0000000;
		Dplus[2583] = 14'b0000000_0000000;
		Dplus[2584] = 14'b0000000_0000000;
		Dplus[2585] = 14'b0000000_0000000;
		Dplus[2586] = 14'b0000000_0000000;
		Dplus[2587] = 14'b0000000_0000000;
		Dplus[2588] = 14'b0000000_0000000;
		Dplus[2589] = 14'b0000000_0000000;
		Dplus[2590] = 14'b0000000_0000000;
		Dplus[2591] = 14'b0000000_0000000;
		Dplus[2592] = 14'b0000000_0000000;
		Dplus[2593] = 14'b0000000_0000000;
		Dplus[2594] = 14'b0000000_0000000;
		Dplus[2595] = 14'b0000000_0000000;
		Dplus[2596] = 14'b0000000_0000000;
		Dplus[2597] = 14'b0000000_0000000;
		Dplus[2598] = 14'b0000000_0000000;
		Dplus[2599] = 14'b0000000_0000000;
		Dplus[2600] = 14'b0000000_0000000;
		Dplus[2601] = 14'b0000000_0000000;
		Dplus[2602] = 14'b0000000_0000000;
		Dplus[2603] = 14'b0000000_0000000;
		Dplus[2604] = 14'b0000000_0000000;
		Dplus[2605] = 14'b0000000_0000000;
		Dplus[2606] = 14'b0000000_0000000;
		Dplus[2607] = 14'b0000000_0000000;
		Dplus[2608] = 14'b0000000_0000000;
		Dplus[2609] = 14'b0000000_0000000;
		Dplus[2610] = 14'b0000000_0000000;
		Dplus[2611] = 14'b0000000_0000000;
		Dplus[2612] = 14'b0000000_0000000;
		Dplus[2613] = 14'b0000000_0000000;
		Dplus[2614] = 14'b0000000_0000000;
		Dplus[2615] = 14'b0000000_0000000;
		Dplus[2616] = 14'b0000000_0000000;
		Dplus[2617] = 14'b0000000_0000000;
		Dplus[2618] = 14'b0000000_0000000;
		Dplus[2619] = 14'b0000000_0000000;
		Dplus[2620] = 14'b0000000_0000000;
		Dplus[2621] = 14'b0000000_0000000;
		Dplus[2622] = 14'b0000000_0000000;
		Dplus[2623] = 14'b0000000_0000000;
		Dplus[2624] = 14'b0000000_0000000;
		Dplus[2625] = 14'b0000000_0000000;
		Dplus[2626] = 14'b0000000_0000000;
		Dplus[2627] = 14'b0000000_0000000;
		Dplus[2628] = 14'b0000000_0000000;
		Dplus[2629] = 14'b0000000_0000000;
		Dplus[2630] = 14'b0000000_0000000;
		Dplus[2631] = 14'b0000000_0000000;
		Dplus[2632] = 14'b0000000_0000000;
		Dplus[2633] = 14'b0000000_0000000;
		Dplus[2634] = 14'b0000000_0000000;
		Dplus[2635] = 14'b0000000_0000000;
		Dplus[2636] = 14'b0000000_0000000;
		Dplus[2637] = 14'b0000000_0000000;
		Dplus[2638] = 14'b0000000_0000000;
		Dplus[2639] = 14'b0000000_0000000;
		Dplus[2640] = 14'b0000000_0000000;
		Dplus[2641] = 14'b0000000_0000000;
		Dplus[2642] = 14'b0000000_0000000;
		Dplus[2643] = 14'b0000000_0000000;
		Dplus[2644] = 14'b0000000_0000000;
		Dplus[2645] = 14'b0000000_0000000;
		Dplus[2646] = 14'b0000000_0000000;
		Dplus[2647] = 14'b0000000_0000000;
		Dplus[2648] = 14'b0000000_0000000;
		Dplus[2649] = 14'b0000000_0000000;
		Dplus[2650] = 14'b0000000_0000000;
		Dplus[2651] = 14'b0000000_0000000;
		Dplus[2652] = 14'b0000000_0000000;
		Dplus[2653] = 14'b0000000_0000000;
		Dplus[2654] = 14'b0000000_0000000;
		Dplus[2655] = 14'b0000000_0000000;
		Dplus[2656] = 14'b0000000_0000000;
		Dplus[2657] = 14'b0000000_0000000;
		Dplus[2658] = 14'b0000000_0000000;
		Dplus[2659] = 14'b0000000_0000000;
		Dplus[2660] = 14'b0000000_0000000;
		Dplus[2661] = 14'b0000000_0000000;
		Dplus[2662] = 14'b0000000_0000000;
		Dplus[2663] = 14'b0000000_0000000;
		Dplus[2664] = 14'b0000000_0000000;
		Dplus[2665] = 14'b0000000_0000000;
		Dplus[2666] = 14'b0000000_0000000;
		Dplus[2667] = 14'b0000000_0000000;
		Dplus[2668] = 14'b0000000_0000000;
		Dplus[2669] = 14'b0000000_0000000;
		Dplus[2670] = 14'b0000000_0000000;
		Dplus[2671] = 14'b0000000_0000000;
		Dplus[2672] = 14'b0000000_0000000;
		Dplus[2673] = 14'b0000000_0000000;
		Dplus[2674] = 14'b0000000_0000000;
		Dplus[2675] = 14'b0000000_0000000;
		Dplus[2676] = 14'b0000000_0000000;
		Dplus[2677] = 14'b0000000_0000000;
		Dplus[2678] = 14'b0000000_0000000;
		Dplus[2679] = 14'b0000000_0000000;
		Dplus[2680] = 14'b0000000_0000000;
		Dplus[2681] = 14'b0000000_0000000;
		Dplus[2682] = 14'b0000000_0000000;
		Dplus[2683] = 14'b0000000_0000000;
		Dplus[2684] = 14'b0000000_0000000;
		Dplus[2685] = 14'b0000000_0000000;
		Dplus[2686] = 14'b0000000_0000000;
		Dplus[2687] = 14'b0000000_0000000;
		Dplus[2688] = 14'b0000000_0000000;
		Dplus[2689] = 14'b0000000_0000000;
		Dplus[2690] = 14'b0000000_0000000;
		Dplus[2691] = 14'b0000000_0000000;
		Dplus[2692] = 14'b0000000_0000000;
		Dplus[2693] = 14'b0000000_0000000;
		Dplus[2694] = 14'b0000000_0000000;
		Dplus[2695] = 14'b0000000_0000000;
		Dplus[2696] = 14'b0000000_0000000;
		Dplus[2697] = 14'b0000000_0000000;
		Dplus[2698] = 14'b0000000_0000000;
		Dplus[2699] = 14'b0000000_0000000;
		Dplus[2700] = 14'b0000000_0000000;
		Dplus[2701] = 14'b0000000_0000000;
		Dplus[2702] = 14'b0000000_0000000;
		Dplus[2703] = 14'b0000000_0000000;
		Dplus[2704] = 14'b0000000_0000000;
		Dplus[2705] = 14'b0000000_0000000;
		Dplus[2706] = 14'b0000000_0000000;
		Dplus[2707] = 14'b0000000_0000000;
		Dplus[2708] = 14'b0000000_0000000;
		Dplus[2709] = 14'b0000000_0000000;
		Dplus[2710] = 14'b0000000_0000000;
		Dplus[2711] = 14'b0000000_0000000;
		Dplus[2712] = 14'b0000000_0000000;
		Dplus[2713] = 14'b0000000_0000000;
		Dplus[2714] = 14'b0000000_0000000;
		Dplus[2715] = 14'b0000000_0000000;
		Dplus[2716] = 14'b0000000_0000000;
		Dplus[2717] = 14'b0000000_0000000;
		Dplus[2718] = 14'b0000000_0000000;
		Dplus[2719] = 14'b0000000_0000000;
		Dplus[2720] = 14'b0000000_0000000;
		Dplus[2721] = 14'b0000000_0000000;
		Dplus[2722] = 14'b0000000_0000000;
		Dplus[2723] = 14'b0000000_0000000;
		Dplus[2724] = 14'b0000000_0000000;
		Dplus[2725] = 14'b0000000_0000000;
		Dplus[2726] = 14'b0000000_0000000;
		Dplus[2727] = 14'b0000000_0000000;
		Dplus[2728] = 14'b0000000_0000000;
		Dplus[2729] = 14'b0000000_0000000;
		Dplus[2730] = 14'b0000000_0000000;
		Dplus[2731] = 14'b0000000_0000000;
		Dplus[2732] = 14'b0000000_0000000;
		Dplus[2733] = 14'b0000000_0000000;
		Dplus[2734] = 14'b0000000_0000000;
		Dplus[2735] = 14'b0000000_0000000;
		Dplus[2736] = 14'b0000000_0000000;
		Dplus[2737] = 14'b0000000_0000000;
		Dplus[2738] = 14'b0000000_0000000;
		Dplus[2739] = 14'b0000000_0000000;
		Dplus[2740] = 14'b0000000_0000000;
		Dplus[2741] = 14'b0000000_0000000;
		Dplus[2742] = 14'b0000000_0000000;
		Dplus[2743] = 14'b0000000_0000000;
		Dplus[2744] = 14'b0000000_0000000;
		Dplus[2745] = 14'b0000000_0000000;
		Dplus[2746] = 14'b0000000_0000000;
		Dplus[2747] = 14'b0000000_0000000;
		Dplus[2748] = 14'b0000000_0000000;
		Dplus[2749] = 14'b0000000_0000000;
		Dplus[2750] = 14'b0000000_0000000;
		Dplus[2751] = 14'b0000000_0000000;
		Dplus[2752] = 14'b0000000_0000000;
		Dplus[2753] = 14'b0000000_0000000;
		Dplus[2754] = 14'b0000000_0000000;
		Dplus[2755] = 14'b0000000_0000000;
		Dplus[2756] = 14'b0000000_0000000;
		Dplus[2757] = 14'b0000000_0000000;
		Dplus[2758] = 14'b0000000_0000000;
		Dplus[2759] = 14'b0000000_0000000;
		Dplus[2760] = 14'b0000000_0000000;
		Dplus[2761] = 14'b0000000_0000000;
		Dplus[2762] = 14'b0000000_0000000;
		Dplus[2763] = 14'b0000000_0000000;
		Dplus[2764] = 14'b0000000_0000000;
		Dplus[2765] = 14'b0000000_0000000;
		Dplus[2766] = 14'b0000000_0000000;
		Dplus[2767] = 14'b0000000_0000000;
		Dplus[2768] = 14'b0000000_0000000;
		Dplus[2769] = 14'b0000000_0000000;
		Dplus[2770] = 14'b0000000_0000000;
		Dplus[2771] = 14'b0000000_0000000;
		Dplus[2772] = 14'b0000000_0000000;
		Dplus[2773] = 14'b0000000_0000000;
		Dplus[2774] = 14'b0000000_0000000;
		Dplus[2775] = 14'b0000000_0000000;
		Dplus[2776] = 14'b0000000_0000000;
		Dplus[2777] = 14'b0000000_0000000;
		Dplus[2778] = 14'b0000000_0000000;
		Dplus[2779] = 14'b0000000_0000000;
		Dplus[2780] = 14'b0000000_0000000;
		Dplus[2781] = 14'b0000000_0000000;
		Dplus[2782] = 14'b0000000_0000000;
		Dplus[2783] = 14'b0000000_0000000;
		Dplus[2784] = 14'b0000000_0000000;
		Dplus[2785] = 14'b0000000_0000000;
		Dplus[2786] = 14'b0000000_0000000;
		Dplus[2787] = 14'b0000000_0000000;
		Dplus[2788] = 14'b0000000_0000000;
		Dplus[2789] = 14'b0000000_0000000;
		Dplus[2790] = 14'b0000000_0000000;
		Dplus[2791] = 14'b0000000_0000000;
		Dplus[2792] = 14'b0000000_0000000;
		Dplus[2793] = 14'b0000000_0000000;
		Dplus[2794] = 14'b0000000_0000000;
		Dplus[2795] = 14'b0000000_0000000;
		Dplus[2796] = 14'b0000000_0000000;
		Dplus[2797] = 14'b0000000_0000000;
		Dplus[2798] = 14'b0000000_0000000;
		Dplus[2799] = 14'b0000000_0000000;
		Dplus[2800] = 14'b0000000_0000000;
		Dplus[2801] = 14'b0000000_0000000;
		Dplus[2802] = 14'b0000000_0000000;
		Dplus[2803] = 14'b0000000_0000000;
		Dplus[2804] = 14'b0000000_0000000;
		Dplus[2805] = 14'b0000000_0000000;
		Dplus[2806] = 14'b0000000_0000000;
		Dplus[2807] = 14'b0000000_0000000;
		Dplus[2808] = 14'b0000000_0000000;
		Dplus[2809] = 14'b0000000_0000000;
		Dplus[2810] = 14'b0000000_0000000;
		Dplus[2811] = 14'b0000000_0000000;
		Dplus[2812] = 14'b0000000_0000000;
		Dplus[2813] = 14'b0000000_0000000;
		Dplus[2814] = 14'b0000000_0000000;
		Dplus[2815] = 14'b0000000_0000000;
		Dplus[2816] = 14'b0000000_0000000;
		Dplus[2817] = 14'b0000000_0000000;
		Dplus[2818] = 14'b0000000_0000000;
		Dplus[2819] = 14'b0000000_0000000;
		Dplus[2820] = 14'b0000000_0000000;
		Dplus[2821] = 14'b0000000_0000000;
		Dplus[2822] = 14'b0000000_0000000;
		Dplus[2823] = 14'b0000000_0000000;
		Dplus[2824] = 14'b0000000_0000000;
		Dplus[2825] = 14'b0000000_0000000;
		Dplus[2826] = 14'b0000000_0000000;
		Dplus[2827] = 14'b0000000_0000000;
		Dplus[2828] = 14'b0000000_0000000;
		Dplus[2829] = 14'b0000000_0000000;
		Dplus[2830] = 14'b0000000_0000000;
		Dplus[2831] = 14'b0000000_0000000;
		Dplus[2832] = 14'b0000000_0000000;
		Dplus[2833] = 14'b0000000_0000000;
		Dplus[2834] = 14'b0000000_0000000;
		Dplus[2835] = 14'b0000000_0000000;
		Dplus[2836] = 14'b0000000_0000000;
		Dplus[2837] = 14'b0000000_0000000;
		Dplus[2838] = 14'b0000000_0000000;
		Dplus[2839] = 14'b0000000_0000000;
		Dplus[2840] = 14'b0000000_0000000;
		Dplus[2841] = 14'b0000000_0000000;
		Dplus[2842] = 14'b0000000_0000000;
		Dplus[2843] = 14'b0000000_0000000;
		Dplus[2844] = 14'b0000000_0000000;
		Dplus[2845] = 14'b0000000_0000000;
		Dplus[2846] = 14'b0000000_0000000;
		Dplus[2847] = 14'b0000000_0000000;
		Dplus[2848] = 14'b0000000_0000000;
		Dplus[2849] = 14'b0000000_0000000;
		Dplus[2850] = 14'b0000000_0000000;
		Dplus[2851] = 14'b0000000_0000000;
		Dplus[2852] = 14'b0000000_0000000;
		Dplus[2853] = 14'b0000000_0000000;
		Dplus[2854] = 14'b0000000_0000000;
		Dplus[2855] = 14'b0000000_0000000;
		Dplus[2856] = 14'b0000000_0000000;
		Dplus[2857] = 14'b0000000_0000000;
		Dplus[2858] = 14'b0000000_0000000;
		Dplus[2859] = 14'b0000000_0000000;
		Dplus[2860] = 14'b0000000_0000000;
		Dplus[2861] = 14'b0000000_0000000;
		Dplus[2862] = 14'b0000000_0000000;
		Dplus[2863] = 14'b0000000_0000000;
		Dplus[2864] = 14'b0000000_0000000;
		Dplus[2865] = 14'b0000000_0000000;
		Dplus[2866] = 14'b0000000_0000000;
		Dplus[2867] = 14'b0000000_0000000;
		Dplus[2868] = 14'b0000000_0000000;
		Dplus[2869] = 14'b0000000_0000000;
		Dplus[2870] = 14'b0000000_0000000;
		Dplus[2871] = 14'b0000000_0000000;
		Dplus[2872] = 14'b0000000_0000000;
		Dplus[2873] = 14'b0000000_0000000;
		Dplus[2874] = 14'b0000000_0000000;
		Dplus[2875] = 14'b0000000_0000000;
		Dplus[2876] = 14'b0000000_0000000;
		Dplus[2877] = 14'b0000000_0000000;
		Dplus[2878] = 14'b0000000_0000000;
		Dplus[2879] = 14'b0000000_0000000;
		Dplus[2880] = 14'b0000000_0000000;
		Dplus[2881] = 14'b0000000_0000000;
		Dplus[2882] = 14'b0000000_0000000;
		Dplus[2883] = 14'b0000000_0000000;
		Dplus[2884] = 14'b0000000_0000000;
		Dplus[2885] = 14'b0000000_0000000;
		Dplus[2886] = 14'b0000000_0000000;
		Dplus[2887] = 14'b0000000_0000000;
		Dplus[2888] = 14'b0000000_0000000;
		Dplus[2889] = 14'b0000000_0000000;
		Dplus[2890] = 14'b0000000_0000000;
		Dplus[2891] = 14'b0000000_0000000;
		Dplus[2892] = 14'b0000000_0000000;
		Dplus[2893] = 14'b0000000_0000000;
		Dplus[2894] = 14'b0000000_0000000;
		Dplus[2895] = 14'b0000000_0000000;
		Dplus[2896] = 14'b0000000_0000000;
		Dplus[2897] = 14'b0000000_0000000;
		Dplus[2898] = 14'b0000000_0000000;
		Dplus[2899] = 14'b0000000_0000000;
		Dplus[2900] = 14'b0000000_0000000;
		Dplus[2901] = 14'b0000000_0000000;
		Dplus[2902] = 14'b0000000_0000000;
		Dplus[2903] = 14'b0000000_0000000;
		Dplus[2904] = 14'b0000000_0000000;
		Dplus[2905] = 14'b0000000_0000000;
		Dplus[2906] = 14'b0000000_0000000;
		Dplus[2907] = 14'b0000000_0000000;
		Dplus[2908] = 14'b0000000_0000000;
		Dplus[2909] = 14'b0000000_0000000;
		Dplus[2910] = 14'b0000000_0000000;
		Dplus[2911] = 14'b0000000_0000000;
		Dplus[2912] = 14'b0000000_0000000;
		Dplus[2913] = 14'b0000000_0000000;
		Dplus[2914] = 14'b0000000_0000000;
		Dplus[2915] = 14'b0000000_0000000;
		Dplus[2916] = 14'b0000000_0000000;
		Dplus[2917] = 14'b0000000_0000000;
		Dplus[2918] = 14'b0000000_0000000;
		Dplus[2919] = 14'b0000000_0000000;
		Dplus[2920] = 14'b0000000_0000000;
		Dplus[2921] = 14'b0000000_0000000;
		Dplus[2922] = 14'b0000000_0000000;
		Dplus[2923] = 14'b0000000_0000000;
		Dplus[2924] = 14'b0000000_0000000;
		Dplus[2925] = 14'b0000000_0000000;
		Dplus[2926] = 14'b0000000_0000000;
		Dplus[2927] = 14'b0000000_0000000;
		Dplus[2928] = 14'b0000000_0000000;
		Dplus[2929] = 14'b0000000_0000000;
		Dplus[2930] = 14'b0000000_0000000;
		Dplus[2931] = 14'b0000000_0000000;
		Dplus[2932] = 14'b0000000_0000000;
		Dplus[2933] = 14'b0000000_0000000;
		Dplus[2934] = 14'b0000000_0000000;
		Dplus[2935] = 14'b0000000_0000000;
		Dplus[2936] = 14'b0000000_0000000;
		Dplus[2937] = 14'b0000000_0000000;
		Dplus[2938] = 14'b0000000_0000000;
		Dplus[2939] = 14'b0000000_0000000;
		Dplus[2940] = 14'b0000000_0000000;
		Dplus[2941] = 14'b0000000_0000000;
		Dplus[2942] = 14'b0000000_0000000;
		Dplus[2943] = 14'b0000000_0000000;
		Dplus[2944] = 14'b0000000_0000000;
		Dplus[2945] = 14'b0000000_0000000;
		Dplus[2946] = 14'b0000000_0000000;
		Dplus[2947] = 14'b0000000_0000000;
		Dplus[2948] = 14'b0000000_0000000;
		Dplus[2949] = 14'b0000000_0000000;
		Dplus[2950] = 14'b0000000_0000000;
		Dplus[2951] = 14'b0000000_0000000;
		Dplus[2952] = 14'b0000000_0000000;
		Dplus[2953] = 14'b0000000_0000000;
		Dplus[2954] = 14'b0000000_0000000;
		Dplus[2955] = 14'b0000000_0000000;
		Dplus[2956] = 14'b0000000_0000000;
		Dplus[2957] = 14'b0000000_0000000;
		Dplus[2958] = 14'b0000000_0000000;
		Dplus[2959] = 14'b0000000_0000000;
		Dplus[2960] = 14'b0000000_0000000;
		Dplus[2961] = 14'b0000000_0000000;
		Dplus[2962] = 14'b0000000_0000000;
		Dplus[2963] = 14'b0000000_0000000;
		Dplus[2964] = 14'b0000000_0000000;
		Dplus[2965] = 14'b0000000_0000000;
		Dplus[2966] = 14'b0000000_0000000;
		Dplus[2967] = 14'b0000000_0000000;
		Dplus[2968] = 14'b0000000_0000000;
		Dplus[2969] = 14'b0000000_0000000;
		Dplus[2970] = 14'b0000000_0000000;
		Dplus[2971] = 14'b0000000_0000000;
		Dplus[2972] = 14'b0000000_0000000;
		Dplus[2973] = 14'b0000000_0000000;
		Dplus[2974] = 14'b0000000_0000000;
		Dplus[2975] = 14'b0000000_0000000;
		Dplus[2976] = 14'b0000000_0000000;
		Dplus[2977] = 14'b0000000_0000000;
		Dplus[2978] = 14'b0000000_0000000;
		Dplus[2979] = 14'b0000000_0000000;
		Dplus[2980] = 14'b0000000_0000000;
		Dplus[2981] = 14'b0000000_0000000;
		Dplus[2982] = 14'b0000000_0000000;
		Dplus[2983] = 14'b0000000_0000000;
		Dplus[2984] = 14'b0000000_0000000;
		Dplus[2985] = 14'b0000000_0000000;
		Dplus[2986] = 14'b0000000_0000000;
		Dplus[2987] = 14'b0000000_0000000;
		Dplus[2988] = 14'b0000000_0000000;
		Dplus[2989] = 14'b0000000_0000000;
		Dplus[2990] = 14'b0000000_0000000;
		Dplus[2991] = 14'b0000000_0000000;
		Dplus[2992] = 14'b0000000_0000000;
		Dplus[2993] = 14'b0000000_0000000;
		Dplus[2994] = 14'b0000000_0000000;
		Dplus[2995] = 14'b0000000_0000000;
		Dplus[2996] = 14'b0000000_0000000;
		Dplus[2997] = 14'b0000000_0000000;
		Dplus[2998] = 14'b0000000_0000000;
		Dplus[2999] = 14'b0000000_0000000;
		Dplus[3000] = 14'b0000000_0000000;
		Dplus[3001] = 14'b0000000_0000000;
		Dplus[3002] = 14'b0000000_0000000;
		Dplus[3003] = 14'b0000000_0000000;
		Dplus[3004] = 14'b0000000_0000000;
		Dplus[3005] = 14'b0000000_0000000;
		Dplus[3006] = 14'b0000000_0000000;
		Dplus[3007] = 14'b0000000_0000000;
		Dplus[3008] = 14'b0000000_0000000;
		Dplus[3009] = 14'b0000000_0000000;
		Dplus[3010] = 14'b0000000_0000000;
		Dplus[3011] = 14'b0000000_0000000;
		Dplus[3012] = 14'b0000000_0000000;
		Dplus[3013] = 14'b0000000_0000000;
		Dplus[3014] = 14'b0000000_0000000;
		Dplus[3015] = 14'b0000000_0000000;
		Dplus[3016] = 14'b0000000_0000000;
		Dplus[3017] = 14'b0000000_0000000;
		Dplus[3018] = 14'b0000000_0000000;
		Dplus[3019] = 14'b0000000_0000000;
		Dplus[3020] = 14'b0000000_0000000;
		Dplus[3021] = 14'b0000000_0000000;
		Dplus[3022] = 14'b0000000_0000000;
		Dplus[3023] = 14'b0000000_0000000;
		Dplus[3024] = 14'b0000000_0000000;
		Dplus[3025] = 14'b0000000_0000000;
		Dplus[3026] = 14'b0000000_0000000;
		Dplus[3027] = 14'b0000000_0000000;
		Dplus[3028] = 14'b0000000_0000000;
		Dplus[3029] = 14'b0000000_0000000;
		Dplus[3030] = 14'b0000000_0000000;
		Dplus[3031] = 14'b0000000_0000000;
		Dplus[3032] = 14'b0000000_0000000;
		Dplus[3033] = 14'b0000000_0000000;
		Dplus[3034] = 14'b0000000_0000000;
		Dplus[3035] = 14'b0000000_0000000;
		Dplus[3036] = 14'b0000000_0000000;
		Dplus[3037] = 14'b0000000_0000000;
		Dplus[3038] = 14'b0000000_0000000;
		Dplus[3039] = 14'b0000000_0000000;
		Dplus[3040] = 14'b0000000_0000000;
		Dplus[3041] = 14'b0000000_0000000;
		Dplus[3042] = 14'b0000000_0000000;
		Dplus[3043] = 14'b0000000_0000000;
		Dplus[3044] = 14'b0000000_0000000;
		Dplus[3045] = 14'b0000000_0000000;
		Dplus[3046] = 14'b0000000_0000000;
		Dplus[3047] = 14'b0000000_0000000;
		Dplus[3048] = 14'b0000000_0000000;
		Dplus[3049] = 14'b0000000_0000000;
		Dplus[3050] = 14'b0000000_0000000;
		Dplus[3051] = 14'b0000000_0000000;
		Dplus[3052] = 14'b0000000_0000000;
		Dplus[3053] = 14'b0000000_0000000;
		Dplus[3054] = 14'b0000000_0000000;
		Dplus[3055] = 14'b0000000_0000000;
		Dplus[3056] = 14'b0000000_0000000;
		Dplus[3057] = 14'b0000000_0000000;
		Dplus[3058] = 14'b0000000_0000000;
		Dplus[3059] = 14'b0000000_0000000;
		Dplus[3060] = 14'b0000000_0000000;
		Dplus[3061] = 14'b0000000_0000000;
		Dplus[3062] = 14'b0000000_0000000;
		Dplus[3063] = 14'b0000000_0000000;
		Dplus[3064] = 14'b0000000_0000000;
		Dplus[3065] = 14'b0000000_0000000;
		Dplus[3066] = 14'b0000000_0000000;
		Dplus[3067] = 14'b0000000_0000000;
		Dplus[3068] = 14'b0000000_0000000;
		Dplus[3069] = 14'b0000000_0000000;
		Dplus[3070] = 14'b0000000_0000000;
		Dplus[3071] = 14'b0000000_0000000;
		Dplus[3072] = 14'b0000000_0000000;
		Dplus[3073] = 14'b0000000_0000000;
		Dplus[3074] = 14'b0000000_0000000;
		Dplus[3075] = 14'b0000000_0000000;
		Dplus[3076] = 14'b0000000_0000000;
		Dplus[3077] = 14'b0000000_0000000;
		Dplus[3078] = 14'b0000000_0000000;
		Dplus[3079] = 14'b0000000_0000000;
		Dplus[3080] = 14'b0000000_0000000;
		Dplus[3081] = 14'b0000000_0000000;
		Dplus[3082] = 14'b0000000_0000000;
		Dplus[3083] = 14'b0000000_0000000;
		Dplus[3084] = 14'b0000000_0000000;
		Dplus[3085] = 14'b0000000_0000000;
		Dplus[3086] = 14'b0000000_0000000;
		Dplus[3087] = 14'b0000000_0000000;
		Dplus[3088] = 14'b0000000_0000000;
		Dplus[3089] = 14'b0000000_0000000;
		Dplus[3090] = 14'b0000000_0000000;
		Dplus[3091] = 14'b0000000_0000000;
		Dplus[3092] = 14'b0000000_0000000;
		Dplus[3093] = 14'b0000000_0000000;
		Dplus[3094] = 14'b0000000_0000000;
		Dplus[3095] = 14'b0000000_0000000;
		Dplus[3096] = 14'b0000000_0000000;
		Dplus[3097] = 14'b0000000_0000000;
		Dplus[3098] = 14'b0000000_0000000;
		Dplus[3099] = 14'b0000000_0000000;
		Dplus[3100] = 14'b0000000_0000000;
		Dplus[3101] = 14'b0000000_0000000;
		Dplus[3102] = 14'b0000000_0000000;
		Dplus[3103] = 14'b0000000_0000000;
		Dplus[3104] = 14'b0000000_0000000;
		Dplus[3105] = 14'b0000000_0000000;
		Dplus[3106] = 14'b0000000_0000000;
		Dplus[3107] = 14'b0000000_0000000;
		Dplus[3108] = 14'b0000000_0000000;
		Dplus[3109] = 14'b0000000_0000000;
		Dplus[3110] = 14'b0000000_0000000;
		Dplus[3111] = 14'b0000000_0000000;
		Dplus[3112] = 14'b0000000_0000000;
		Dplus[3113] = 14'b0000000_0000000;
		Dplus[3114] = 14'b0000000_0000000;
		Dplus[3115] = 14'b0000000_0000000;
		Dplus[3116] = 14'b0000000_0000000;
		Dplus[3117] = 14'b0000000_0000000;
		Dplus[3118] = 14'b0000000_0000000;
		Dplus[3119] = 14'b0000000_0000000;
		Dplus[3120] = 14'b0000000_0000000;
		Dplus[3121] = 14'b0000000_0000000;
		Dplus[3122] = 14'b0000000_0000000;
		Dplus[3123] = 14'b0000000_0000000;
		Dplus[3124] = 14'b0000000_0000000;
		Dplus[3125] = 14'b0000000_0000000;
		Dplus[3126] = 14'b0000000_0000000;
		Dplus[3127] = 14'b0000000_0000000;
		Dplus[3128] = 14'b0000000_0000000;
		Dplus[3129] = 14'b0000000_0000000;
		Dplus[3130] = 14'b0000000_0000000;
		Dplus[3131] = 14'b0000000_0000000;
		Dplus[3132] = 14'b0000000_0000000;
		Dplus[3133] = 14'b0000000_0000000;
		Dplus[3134] = 14'b0000000_0000000;
		Dplus[3135] = 14'b0000000_0000000;
		Dplus[3136] = 14'b0000000_0000000;
		Dplus[3137] = 14'b0000000_0000000;
		Dplus[3138] = 14'b0000000_0000000;
		Dplus[3139] = 14'b0000000_0000000;
		Dplus[3140] = 14'b0000000_0000000;
		Dplus[3141] = 14'b0000000_0000000;
		Dplus[3142] = 14'b0000000_0000000;
		Dplus[3143] = 14'b0000000_0000000;
		Dplus[3144] = 14'b0000000_0000000;
		Dplus[3145] = 14'b0000000_0000000;
		Dplus[3146] = 14'b0000000_0000000;
		Dplus[3147] = 14'b0000000_0000000;
		Dplus[3148] = 14'b0000000_0000000;
		Dplus[3149] = 14'b0000000_0000000;
		Dplus[3150] = 14'b0000000_0000000;
		Dplus[3151] = 14'b0000000_0000000;
		Dplus[3152] = 14'b0000000_0000000;
		Dplus[3153] = 14'b0000000_0000000;
		Dplus[3154] = 14'b0000000_0000000;
		Dplus[3155] = 14'b0000000_0000000;
		Dplus[3156] = 14'b0000000_0000000;
		Dplus[3157] = 14'b0000000_0000000;
		Dplus[3158] = 14'b0000000_0000000;
		Dplus[3159] = 14'b0000000_0000000;
		Dplus[3160] = 14'b0000000_0000000;
		Dplus[3161] = 14'b0000000_0000000;
		Dplus[3162] = 14'b0000000_0000000;
		Dplus[3163] = 14'b0000000_0000000;
		Dplus[3164] = 14'b0000000_0000000;
		Dplus[3165] = 14'b0000000_0000000;
		Dplus[3166] = 14'b0000000_0000000;
		Dplus[3167] = 14'b0000000_0000000;
		Dplus[3168] = 14'b0000000_0000000;
		Dplus[3169] = 14'b0000000_0000000;
		Dplus[3170] = 14'b0000000_0000000;
		Dplus[3171] = 14'b0000000_0000000;
		Dplus[3172] = 14'b0000000_0000000;
		Dplus[3173] = 14'b0000000_0000000;
		Dplus[3174] = 14'b0000000_0000000;
		Dplus[3175] = 14'b0000000_0000000;
		Dplus[3176] = 14'b0000000_0000000;
		Dplus[3177] = 14'b0000000_0000000;
		Dplus[3178] = 14'b0000000_0000000;
		Dplus[3179] = 14'b0000000_0000000;
		Dplus[3180] = 14'b0000000_0000000;
		Dplus[3181] = 14'b0000000_0000000;
		Dplus[3182] = 14'b0000000_0000000;
		Dplus[3183] = 14'b0000000_0000000;
		Dplus[3184] = 14'b0000000_0000000;
		Dplus[3185] = 14'b0000000_0000000;
		Dplus[3186] = 14'b0000000_0000000;
		Dplus[3187] = 14'b0000000_0000000;
		Dplus[3188] = 14'b0000000_0000000;
		Dplus[3189] = 14'b0000000_0000000;
		Dplus[3190] = 14'b0000000_0000000;
		Dplus[3191] = 14'b0000000_0000000;
		Dplus[3192] = 14'b0000000_0000000;
		Dplus[3193] = 14'b0000000_0000000;
		Dplus[3194] = 14'b0000000_0000000;
		Dplus[3195] = 14'b0000000_0000000;
		Dplus[3196] = 14'b0000000_0000000;
		Dplus[3197] = 14'b0000000_0000000;
		Dplus[3198] = 14'b0000000_0000000;
		Dplus[3199] = 14'b0000000_0000000;
		Dplus[3200] = 14'b0000000_0000000;
		Dplus[3201] = 14'b0000000_0000000;
		Dplus[3202] = 14'b0000000_0000000;
		Dplus[3203] = 14'b0000000_0000000;
		Dplus[3204] = 14'b0000000_0000000;
		Dplus[3205] = 14'b0000000_0000000;
		Dplus[3206] = 14'b0000000_0000000;
		Dplus[3207] = 14'b0000000_0000000;
		Dplus[3208] = 14'b0000000_0000000;
		Dplus[3209] = 14'b0000000_0000000;
		Dplus[3210] = 14'b0000000_0000000;
		Dplus[3211] = 14'b0000000_0000000;
		Dplus[3212] = 14'b0000000_0000000;
		Dplus[3213] = 14'b0000000_0000000;
		Dplus[3214] = 14'b0000000_0000000;
		Dplus[3215] = 14'b0000000_0000000;
		Dplus[3216] = 14'b0000000_0000000;
		Dplus[3217] = 14'b0000000_0000000;
		Dplus[3218] = 14'b0000000_0000000;
		Dplus[3219] = 14'b0000000_0000000;
		Dplus[3220] = 14'b0000000_0000000;
		Dplus[3221] = 14'b0000000_0000000;
		Dplus[3222] = 14'b0000000_0000000;
		Dplus[3223] = 14'b0000000_0000000;
		Dplus[3224] = 14'b0000000_0000000;
		Dplus[3225] = 14'b0000000_0000000;
		Dplus[3226] = 14'b0000000_0000000;
		Dplus[3227] = 14'b0000000_0000000;
		Dplus[3228] = 14'b0000000_0000000;
		Dplus[3229] = 14'b0000000_0000000;
		Dplus[3230] = 14'b0000000_0000000;
		Dplus[3231] = 14'b0000000_0000000;
		Dplus[3232] = 14'b0000000_0000000;
		Dplus[3233] = 14'b0000000_0000000;
		Dplus[3234] = 14'b0000000_0000000;
		Dplus[3235] = 14'b0000000_0000000;
		Dplus[3236] = 14'b0000000_0000000;
		Dplus[3237] = 14'b0000000_0000000;
		Dplus[3238] = 14'b0000000_0000000;
		Dplus[3239] = 14'b0000000_0000000;
		Dplus[3240] = 14'b0000000_0000000;
		Dplus[3241] = 14'b0000000_0000000;
		Dplus[3242] = 14'b0000000_0000000;
		Dplus[3243] = 14'b0000000_0000000;
		Dplus[3244] = 14'b0000000_0000000;
		Dplus[3245] = 14'b0000000_0000000;
		Dplus[3246] = 14'b0000000_0000000;
		Dplus[3247] = 14'b0000000_0000000;
		Dplus[3248] = 14'b0000000_0000000;
		Dplus[3249] = 14'b0000000_0000000;
		Dplus[3250] = 14'b0000000_0000000;
		Dplus[3251] = 14'b0000000_0000000;
		Dplus[3252] = 14'b0000000_0000000;
		Dplus[3253] = 14'b0000000_0000000;
		Dplus[3254] = 14'b0000000_0000000;
		Dplus[3255] = 14'b0000000_0000000;
		Dplus[3256] = 14'b0000000_0000000;
		Dplus[3257] = 14'b0000000_0000000;
		Dplus[3258] = 14'b0000000_0000000;
		Dplus[3259] = 14'b0000000_0000000;
		Dplus[3260] = 14'b0000000_0000000;
		Dplus[3261] = 14'b0000000_0000000;
		Dplus[3262] = 14'b0000000_0000000;
		Dplus[3263] = 14'b0000000_0000000;
		Dplus[3264] = 14'b0000000_0000000;
		Dplus[3265] = 14'b0000000_0000000;
		Dplus[3266] = 14'b0000000_0000000;
		Dplus[3267] = 14'b0000000_0000000;
		Dplus[3268] = 14'b0000000_0000000;
		Dplus[3269] = 14'b0000000_0000000;
		Dplus[3270] = 14'b0000000_0000000;
		Dplus[3271] = 14'b0000000_0000000;
		Dplus[3272] = 14'b0000000_0000000;
		Dplus[3273] = 14'b0000000_0000000;
		Dplus[3274] = 14'b0000000_0000000;
		Dplus[3275] = 14'b0000000_0000000;
		Dplus[3276] = 14'b0000000_0000000;
		Dplus[3277] = 14'b0000000_0000000;
		Dplus[3278] = 14'b0000000_0000000;
		Dplus[3279] = 14'b0000000_0000000;
		Dplus[3280] = 14'b0000000_0000000;
		Dplus[3281] = 14'b0000000_0000000;
		Dplus[3282] = 14'b0000000_0000000;
		Dplus[3283] = 14'b0000000_0000000;
		Dplus[3284] = 14'b0000000_0000000;
		Dplus[3285] = 14'b0000000_0000000;
		Dplus[3286] = 14'b0000000_0000000;
		Dplus[3287] = 14'b0000000_0000000;
		Dplus[3288] = 14'b0000000_0000000;
		Dplus[3289] = 14'b0000000_0000000;
		Dplus[3290] = 14'b0000000_0000000;
		Dplus[3291] = 14'b0000000_0000000;
		Dplus[3292] = 14'b0000000_0000000;
		Dplus[3293] = 14'b0000000_0000000;
		Dplus[3294] = 14'b0000000_0000000;
		Dplus[3295] = 14'b0000000_0000000;
		Dplus[3296] = 14'b0000000_0000000;
		Dplus[3297] = 14'b0000000_0000000;
		Dplus[3298] = 14'b0000000_0000000;
		Dplus[3299] = 14'b0000000_0000000;
		Dplus[3300] = 14'b0000000_0000000;
		Dplus[3301] = 14'b0000000_0000000;
		Dplus[3302] = 14'b0000000_0000000;
		Dplus[3303] = 14'b0000000_0000000;
		Dplus[3304] = 14'b0000000_0000000;
		Dplus[3305] = 14'b0000000_0000000;
		Dplus[3306] = 14'b0000000_0000000;
		Dplus[3307] = 14'b0000000_0000000;
		Dplus[3308] = 14'b0000000_0000000;
		Dplus[3309] = 14'b0000000_0000000;
		Dplus[3310] = 14'b0000000_0000000;
		Dplus[3311] = 14'b0000000_0000000;
		Dplus[3312] = 14'b0000000_0000000;
		Dplus[3313] = 14'b0000000_0000000;
		Dplus[3314] = 14'b0000000_0000000;
		Dplus[3315] = 14'b0000000_0000000;
		Dplus[3316] = 14'b0000000_0000000;
		Dplus[3317] = 14'b0000000_0000000;
		Dplus[3318] = 14'b0000000_0000000;
		Dplus[3319] = 14'b0000000_0000000;
		Dplus[3320] = 14'b0000000_0000000;
		Dplus[3321] = 14'b0000000_0000000;
		Dplus[3322] = 14'b0000000_0000000;
		Dplus[3323] = 14'b0000000_0000000;
		Dplus[3324] = 14'b0000000_0000000;
		Dplus[3325] = 14'b0000000_0000000;
		Dplus[3326] = 14'b0000000_0000000;
		Dplus[3327] = 14'b0000000_0000000;
		Dplus[3328] = 14'b0000000_0000000;
		Dplus[3329] = 14'b0000000_0000000;
		Dplus[3330] = 14'b0000000_0000000;
		Dplus[3331] = 14'b0000000_0000000;
		Dplus[3332] = 14'b0000000_0000000;
		Dplus[3333] = 14'b0000000_0000000;
		Dplus[3334] = 14'b0000000_0000000;
		Dplus[3335] = 14'b0000000_0000000;
		Dplus[3336] = 14'b0000000_0000000;
		Dplus[3337] = 14'b0000000_0000000;
		Dplus[3338] = 14'b0000000_0000000;
		Dplus[3339] = 14'b0000000_0000000;
		Dplus[3340] = 14'b0000000_0000000;
		Dplus[3341] = 14'b0000000_0000000;
		Dplus[3342] = 14'b0000000_0000000;
		Dplus[3343] = 14'b0000000_0000000;
		Dplus[3344] = 14'b0000000_0000000;
		Dplus[3345] = 14'b0000000_0000000;
		Dplus[3346] = 14'b0000000_0000000;
		Dplus[3347] = 14'b0000000_0000000;
		Dplus[3348] = 14'b0000000_0000000;
		Dplus[3349] = 14'b0000000_0000000;
		Dplus[3350] = 14'b0000000_0000000;
		Dplus[3351] = 14'b0000000_0000000;
		Dplus[3352] = 14'b0000000_0000000;
		Dplus[3353] = 14'b0000000_0000000;
		Dplus[3354] = 14'b0000000_0000000;
		Dplus[3355] = 14'b0000000_0000000;
		Dplus[3356] = 14'b0000000_0000000;
		Dplus[3357] = 14'b0000000_0000000;
		Dplus[3358] = 14'b0000000_0000000;
		Dplus[3359] = 14'b0000000_0000000;
		Dplus[3360] = 14'b0000000_0000000;
		Dplus[3361] = 14'b0000000_0000000;
		Dplus[3362] = 14'b0000000_0000000;
		Dplus[3363] = 14'b0000000_0000000;
		Dplus[3364] = 14'b0000000_0000000;
		Dplus[3365] = 14'b0000000_0000000;
		Dplus[3366] = 14'b0000000_0000000;
		Dplus[3367] = 14'b0000000_0000000;
		Dplus[3368] = 14'b0000000_0000000;
		Dplus[3369] = 14'b0000000_0000000;
		Dplus[3370] = 14'b0000000_0000000;
		Dplus[3371] = 14'b0000000_0000000;
		Dplus[3372] = 14'b0000000_0000000;
		Dplus[3373] = 14'b0000000_0000000;
		Dplus[3374] = 14'b0000000_0000000;
		Dplus[3375] = 14'b0000000_0000000;
		Dplus[3376] = 14'b0000000_0000000;
		Dplus[3377] = 14'b0000000_0000000;
		Dplus[3378] = 14'b0000000_0000000;
		Dplus[3379] = 14'b0000000_0000000;
		Dplus[3380] = 14'b0000000_0000000;
		Dplus[3381] = 14'b0000000_0000000;
		Dplus[3382] = 14'b0000000_0000000;
		Dplus[3383] = 14'b0000000_0000000;
		Dplus[3384] = 14'b0000000_0000000;
		Dplus[3385] = 14'b0000000_0000000;
		Dplus[3386] = 14'b0000000_0000000;
		Dplus[3387] = 14'b0000000_0000000;
		Dplus[3388] = 14'b0000000_0000000;
		Dplus[3389] = 14'b0000000_0000000;
		Dplus[3390] = 14'b0000000_0000000;
		Dplus[3391] = 14'b0000000_0000000;
		Dplus[3392] = 14'b0000000_0000000;
		Dplus[3393] = 14'b0000000_0000000;
		Dplus[3394] = 14'b0000000_0000000;
		Dplus[3395] = 14'b0000000_0000000;
		Dplus[3396] = 14'b0000000_0000000;
		Dplus[3397] = 14'b0000000_0000000;
		Dplus[3398] = 14'b0000000_0000000;
		Dplus[3399] = 14'b0000000_0000000;
		Dplus[3400] = 14'b0000000_0000000;
		Dplus[3401] = 14'b0000000_0000000;
		Dplus[3402] = 14'b0000000_0000000;
		Dplus[3403] = 14'b0000000_0000000;
		Dplus[3404] = 14'b0000000_0000000;
		Dplus[3405] = 14'b0000000_0000000;
		Dplus[3406] = 14'b0000000_0000000;
		Dplus[3407] = 14'b0000000_0000000;
		Dplus[3408] = 14'b0000000_0000000;
		Dplus[3409] = 14'b0000000_0000000;
		Dplus[3410] = 14'b0000000_0000000;
		Dplus[3411] = 14'b0000000_0000000;
		Dplus[3412] = 14'b0000000_0000000;
		Dplus[3413] = 14'b0000000_0000000;
		Dplus[3414] = 14'b0000000_0000000;
		Dplus[3415] = 14'b0000000_0000000;
		Dplus[3416] = 14'b0000000_0000000;
		Dplus[3417] = 14'b0000000_0000000;
		Dplus[3418] = 14'b0000000_0000000;
		Dplus[3419] = 14'b0000000_0000000;
		Dplus[3420] = 14'b0000000_0000000;
		Dplus[3421] = 14'b0000000_0000000;
		Dplus[3422] = 14'b0000000_0000000;
		Dplus[3423] = 14'b0000000_0000000;
		Dplus[3424] = 14'b0000000_0000000;
		Dplus[3425] = 14'b0000000_0000000;
		Dplus[3426] = 14'b0000000_0000000;
		Dplus[3427] = 14'b0000000_0000000;
		Dplus[3428] = 14'b0000000_0000000;
		Dplus[3429] = 14'b0000000_0000000;
		Dplus[3430] = 14'b0000000_0000000;
		Dplus[3431] = 14'b0000000_0000000;
		Dplus[3432] = 14'b0000000_0000000;
		Dplus[3433] = 14'b0000000_0000000;
		Dplus[3434] = 14'b0000000_0000000;
		Dplus[3435] = 14'b0000000_0000000;
		Dplus[3436] = 14'b0000000_0000000;
		Dplus[3437] = 14'b0000000_0000000;
		Dplus[3438] = 14'b0000000_0000000;
		Dplus[3439] = 14'b0000000_0000000;
		Dplus[3440] = 14'b0000000_0000000;
		Dplus[3441] = 14'b0000000_0000000;
		Dplus[3442] = 14'b0000000_0000000;
		Dplus[3443] = 14'b0000000_0000000;
		Dplus[3444] = 14'b0000000_0000000;
		Dplus[3445] = 14'b0000000_0000000;
		Dplus[3446] = 14'b0000000_0000000;
		Dplus[3447] = 14'b0000000_0000000;
		Dplus[3448] = 14'b0000000_0000000;
		Dplus[3449] = 14'b0000000_0000000;
		Dplus[3450] = 14'b0000000_0000000;
		Dplus[3451] = 14'b0000000_0000000;
		Dplus[3452] = 14'b0000000_0000000;
		Dplus[3453] = 14'b0000000_0000000;
		Dplus[3454] = 14'b0000000_0000000;
		Dplus[3455] = 14'b0000000_0000000;
		Dplus[3456] = 14'b0000000_0000000;
		Dplus[3457] = 14'b0000000_0000000;
		Dplus[3458] = 14'b0000000_0000000;
		Dplus[3459] = 14'b0000000_0000000;
		Dplus[3460] = 14'b0000000_0000000;
		Dplus[3461] = 14'b0000000_0000000;
		Dplus[3462] = 14'b0000000_0000000;
		Dplus[3463] = 14'b0000000_0000000;
		Dplus[3464] = 14'b0000000_0000000;
		Dplus[3465] = 14'b0000000_0000000;
		Dplus[3466] = 14'b0000000_0000000;
		Dplus[3467] = 14'b0000000_0000000;
		Dplus[3468] = 14'b0000000_0000000;
		Dplus[3469] = 14'b0000000_0000000;
		Dplus[3470] = 14'b0000000_0000000;
		Dplus[3471] = 14'b0000000_0000000;
		Dplus[3472] = 14'b0000000_0000000;
		Dplus[3473] = 14'b0000000_0000000;
		Dplus[3474] = 14'b0000000_0000000;
		Dplus[3475] = 14'b0000000_0000000;
		Dplus[3476] = 14'b0000000_0000000;
		Dplus[3477] = 14'b0000000_0000000;
		Dplus[3478] = 14'b0000000_0000000;
		Dplus[3479] = 14'b0000000_0000000;
		Dplus[3480] = 14'b0000000_0000000;
		Dplus[3481] = 14'b0000000_0000000;
		Dplus[3482] = 14'b0000000_0000000;
		Dplus[3483] = 14'b0000000_0000000;
		Dplus[3484] = 14'b0000000_0000000;
		Dplus[3485] = 14'b0000000_0000000;
		Dplus[3486] = 14'b0000000_0000000;
		Dplus[3487] = 14'b0000000_0000000;
		Dplus[3488] = 14'b0000000_0000000;
		Dplus[3489] = 14'b0000000_0000000;
		Dplus[3490] = 14'b0000000_0000000;
		Dplus[3491] = 14'b0000000_0000000;
		Dplus[3492] = 14'b0000000_0000000;
		Dplus[3493] = 14'b0000000_0000000;
		Dplus[3494] = 14'b0000000_0000000;
		Dplus[3495] = 14'b0000000_0000000;
		Dplus[3496] = 14'b0000000_0000000;
		Dplus[3497] = 14'b0000000_0000000;
		Dplus[3498] = 14'b0000000_0000000;
		Dplus[3499] = 14'b0000000_0000000;
		Dplus[3500] = 14'b0000000_0000000;
		Dplus[3501] = 14'b0000000_0000000;
		Dplus[3502] = 14'b0000000_0000000;
		Dplus[3503] = 14'b0000000_0000000;
		Dplus[3504] = 14'b0000000_0000000;
		Dplus[3505] = 14'b0000000_0000000;
		Dplus[3506] = 14'b0000000_0000000;
		Dplus[3507] = 14'b0000000_0000000;
		Dplus[3508] = 14'b0000000_0000000;
		Dplus[3509] = 14'b0000000_0000000;
		Dplus[3510] = 14'b0000000_0000000;
		Dplus[3511] = 14'b0000000_0000000;
		Dplus[3512] = 14'b0000000_0000000;
		Dplus[3513] = 14'b0000000_0000000;
		Dplus[3514] = 14'b0000000_0000000;
		Dplus[3515] = 14'b0000000_0000000;
		Dplus[3516] = 14'b0000000_0000000;
		Dplus[3517] = 14'b0000000_0000000;
		Dplus[3518] = 14'b0000000_0000000;
		Dplus[3519] = 14'b0000000_0000000;
		Dplus[3520] = 14'b0000000_0000000;
		Dplus[3521] = 14'b0000000_0000000;
		Dplus[3522] = 14'b0000000_0000000;
		Dplus[3523] = 14'b0000000_0000000;
		Dplus[3524] = 14'b0000000_0000000;
		Dplus[3525] = 14'b0000000_0000000;
		Dplus[3526] = 14'b0000000_0000000;
		Dplus[3527] = 14'b0000000_0000000;
		Dplus[3528] = 14'b0000000_0000000;
		Dplus[3529] = 14'b0000000_0000000;
		Dplus[3530] = 14'b0000000_0000000;
		Dplus[3531] = 14'b0000000_0000000;
		Dplus[3532] = 14'b0000000_0000000;
		Dplus[3533] = 14'b0000000_0000000;
		Dplus[3534] = 14'b0000000_0000000;
		Dplus[3535] = 14'b0000000_0000000;
		Dplus[3536] = 14'b0000000_0000000;
		Dplus[3537] = 14'b0000000_0000000;
		Dplus[3538] = 14'b0000000_0000000;
		Dplus[3539] = 14'b0000000_0000000;
		Dplus[3540] = 14'b0000000_0000000;
		Dplus[3541] = 14'b0000000_0000000;
		Dplus[3542] = 14'b0000000_0000000;
		Dplus[3543] = 14'b0000000_0000000;
		Dplus[3544] = 14'b0000000_0000000;
		Dplus[3545] = 14'b0000000_0000000;
		Dplus[3546] = 14'b0000000_0000000;
		Dplus[3547] = 14'b0000000_0000000;
		Dplus[3548] = 14'b0000000_0000000;
		Dplus[3549] = 14'b0000000_0000000;
		Dplus[3550] = 14'b0000000_0000000;
		Dplus[3551] = 14'b0000000_0000000;
		Dplus[3552] = 14'b0000000_0000000;
		Dplus[3553] = 14'b0000000_0000000;
		Dplus[3554] = 14'b0000000_0000000;
		Dplus[3555] = 14'b0000000_0000000;
		Dplus[3556] = 14'b0000000_0000000;
		Dplus[3557] = 14'b0000000_0000000;
		Dplus[3558] = 14'b0000000_0000000;
		Dplus[3559] = 14'b0000000_0000000;
		Dplus[3560] = 14'b0000000_0000000;
		Dplus[3561] = 14'b0000000_0000000;
		Dplus[3562] = 14'b0000000_0000000;
		Dplus[3563] = 14'b0000000_0000000;
		Dplus[3564] = 14'b0000000_0000000;
		Dplus[3565] = 14'b0000000_0000000;
		Dplus[3566] = 14'b0000000_0000000;
		Dplus[3567] = 14'b0000000_0000000;
		Dplus[3568] = 14'b0000000_0000000;
		Dplus[3569] = 14'b0000000_0000000;
		Dplus[3570] = 14'b0000000_0000000;
		Dplus[3571] = 14'b0000000_0000000;
		Dplus[3572] = 14'b0000000_0000000;
		Dplus[3573] = 14'b0000000_0000000;
		Dplus[3574] = 14'b0000000_0000000;
		Dplus[3575] = 14'b0000000_0000000;
		Dplus[3576] = 14'b0000000_0000000;
		Dplus[3577] = 14'b0000000_0000000;
		Dplus[3578] = 14'b0000000_0000000;
		Dplus[3579] = 14'b0000000_0000000;
		Dplus[3580] = 14'b0000000_0000000;
		Dplus[3581] = 14'b0000000_0000000;
		Dplus[3582] = 14'b0000000_0000000;
		Dplus[3583] = 14'b0000000_0000000;
		Dplus[3584] = 14'b0000000_0000000;
		Dplus[3585] = 14'b0000000_0000000;
		Dplus[3586] = 14'b0000000_0000000;
		Dplus[3587] = 14'b0000000_0000000;
		Dplus[3588] = 14'b0000000_0000000;
		Dplus[3589] = 14'b0000000_0000000;
		Dplus[3590] = 14'b0000000_0000000;
		Dplus[3591] = 14'b0000000_0000000;
		Dplus[3592] = 14'b0000000_0000000;
		Dplus[3593] = 14'b0000000_0000000;
		Dplus[3594] = 14'b0000000_0000000;
		Dplus[3595] = 14'b0000000_0000000;
		Dplus[3596] = 14'b0000000_0000000;
		Dplus[3597] = 14'b0000000_0000000;
		Dplus[3598] = 14'b0000000_0000000;
		Dplus[3599] = 14'b0000000_0000000;
		Dplus[3600] = 14'b0000000_0000000;
		Dplus[3601] = 14'b0000000_0000000;
		Dplus[3602] = 14'b0000000_0000000;
		Dplus[3603] = 14'b0000000_0000000;
		Dplus[3604] = 14'b0000000_0000000;
		Dplus[3605] = 14'b0000000_0000000;
		Dplus[3606] = 14'b0000000_0000000;
		Dplus[3607] = 14'b0000000_0000000;
		Dplus[3608] = 14'b0000000_0000000;
		Dplus[3609] = 14'b0000000_0000000;
		Dplus[3610] = 14'b0000000_0000000;
		Dplus[3611] = 14'b0000000_0000000;
		Dplus[3612] = 14'b0000000_0000000;
		Dplus[3613] = 14'b0000000_0000000;
		Dplus[3614] = 14'b0000000_0000000;
		Dplus[3615] = 14'b0000000_0000000;
		Dplus[3616] = 14'b0000000_0000000;
		Dplus[3617] = 14'b0000000_0000000;
		Dplus[3618] = 14'b0000000_0000000;
		Dplus[3619] = 14'b0000000_0000000;
		Dplus[3620] = 14'b0000000_0000000;
		Dplus[3621] = 14'b0000000_0000000;
		Dplus[3622] = 14'b0000000_0000000;
		Dplus[3623] = 14'b0000000_0000000;
		Dplus[3624] = 14'b0000000_0000000;
		Dplus[3625] = 14'b0000000_0000000;
		Dplus[3626] = 14'b0000000_0000000;
		Dplus[3627] = 14'b0000000_0000000;
		Dplus[3628] = 14'b0000000_0000000;
		Dplus[3629] = 14'b0000000_0000000;
		Dplus[3630] = 14'b0000000_0000000;
		Dplus[3631] = 14'b0000000_0000000;
		Dplus[3632] = 14'b0000000_0000000;
		Dplus[3633] = 14'b0000000_0000000;
		Dplus[3634] = 14'b0000000_0000000;
		Dplus[3635] = 14'b0000000_0000000;
		Dplus[3636] = 14'b0000000_0000000;
		Dplus[3637] = 14'b0000000_0000000;
		Dplus[3638] = 14'b0000000_0000000;
		Dplus[3639] = 14'b0000000_0000000;
		Dplus[3640] = 14'b0000000_0000000;
		Dplus[3641] = 14'b0000000_0000000;
		Dplus[3642] = 14'b0000000_0000000;
		Dplus[3643] = 14'b0000000_0000000;
		Dplus[3644] = 14'b0000000_0000000;
		Dplus[3645] = 14'b0000000_0000000;
		Dplus[3646] = 14'b0000000_0000000;
		Dplus[3647] = 14'b0000000_0000000;
		Dplus[3648] = 14'b0000000_0000000;
		Dplus[3649] = 14'b0000000_0000000;
		Dplus[3650] = 14'b0000000_0000000;
		Dplus[3651] = 14'b0000000_0000000;
		Dplus[3652] = 14'b0000000_0000000;
		Dplus[3653] = 14'b0000000_0000000;
		Dplus[3654] = 14'b0000000_0000000;
		Dplus[3655] = 14'b0000000_0000000;
		Dplus[3656] = 14'b0000000_0000000;
		Dplus[3657] = 14'b0000000_0000000;
		Dplus[3658] = 14'b0000000_0000000;
		Dplus[3659] = 14'b0000000_0000000;
		Dplus[3660] = 14'b0000000_0000000;
		Dplus[3661] = 14'b0000000_0000000;
		Dplus[3662] = 14'b0000000_0000000;
		Dplus[3663] = 14'b0000000_0000000;
		Dplus[3664] = 14'b0000000_0000000;
		Dplus[3665] = 14'b0000000_0000000;
		Dplus[3666] = 14'b0000000_0000000;
		Dplus[3667] = 14'b0000000_0000000;
		Dplus[3668] = 14'b0000000_0000000;
		Dplus[3669] = 14'b0000000_0000000;
		Dplus[3670] = 14'b0000000_0000000;
		Dplus[3671] = 14'b0000000_0000000;
		Dplus[3672] = 14'b0000000_0000000;
		Dplus[3673] = 14'b0000000_0000000;
		Dplus[3674] = 14'b0000000_0000000;
		Dplus[3675] = 14'b0000000_0000000;
		Dplus[3676] = 14'b0000000_0000000;
		Dplus[3677] = 14'b0000000_0000000;
		Dplus[3678] = 14'b0000000_0000000;
		Dplus[3679] = 14'b0000000_0000000;
		Dplus[3680] = 14'b0000000_0000000;
		Dplus[3681] = 14'b0000000_0000000;
		Dplus[3682] = 14'b0000000_0000000;
		Dplus[3683] = 14'b0000000_0000000;
		Dplus[3684] = 14'b0000000_0000000;
		Dplus[3685] = 14'b0000000_0000000;
		Dplus[3686] = 14'b0000000_0000000;
		Dplus[3687] = 14'b0000000_0000000;
		Dplus[3688] = 14'b0000000_0000000;
		Dplus[3689] = 14'b0000000_0000000;
		Dplus[3690] = 14'b0000000_0000000;
		Dplus[3691] = 14'b0000000_0000000;
		Dplus[3692] = 14'b0000000_0000000;
		Dplus[3693] = 14'b0000000_0000000;
		Dplus[3694] = 14'b0000000_0000000;
		Dplus[3695] = 14'b0000000_0000000;
		Dplus[3696] = 14'b0000000_0000000;
		Dplus[3697] = 14'b0000000_0000000;
		Dplus[3698] = 14'b0000000_0000000;
		Dplus[3699] = 14'b0000000_0000000;
		Dplus[3700] = 14'b0000000_0000000;
		Dplus[3701] = 14'b0000000_0000000;
		Dplus[3702] = 14'b0000000_0000000;
		Dplus[3703] = 14'b0000000_0000000;
		Dplus[3704] = 14'b0000000_0000000;
		Dplus[3705] = 14'b0000000_0000000;
		Dplus[3706] = 14'b0000000_0000000;
		Dplus[3707] = 14'b0000000_0000000;
		Dplus[3708] = 14'b0000000_0000000;
		Dplus[3709] = 14'b0000000_0000000;
		Dplus[3710] = 14'b0000000_0000000;
		Dplus[3711] = 14'b0000000_0000000;
		Dplus[3712] = 14'b0000000_0000000;
		Dplus[3713] = 14'b0000000_0000000;
		Dplus[3714] = 14'b0000000_0000000;
		Dplus[3715] = 14'b0000000_0000000;
		Dplus[3716] = 14'b0000000_0000000;
		Dplus[3717] = 14'b0000000_0000000;
		Dplus[3718] = 14'b0000000_0000000;
		Dplus[3719] = 14'b0000000_0000000;
		Dplus[3720] = 14'b0000000_0000000;
		Dplus[3721] = 14'b0000000_0000000;
		Dplus[3722] = 14'b0000000_0000000;
		Dplus[3723] = 14'b0000000_0000000;
		Dplus[3724] = 14'b0000000_0000000;
		Dplus[3725] = 14'b0000000_0000000;
		Dplus[3726] = 14'b0000000_0000000;
		Dplus[3727] = 14'b0000000_0000000;
		Dplus[3728] = 14'b0000000_0000000;
		Dplus[3729] = 14'b0000000_0000000;
		Dplus[3730] = 14'b0000000_0000000;
		Dplus[3731] = 14'b0000000_0000000;
		Dplus[3732] = 14'b0000000_0000000;
		Dplus[3733] = 14'b0000000_0000000;
		Dplus[3734] = 14'b0000000_0000000;
		Dplus[3735] = 14'b0000000_0000000;
		Dplus[3736] = 14'b0000000_0000000;
		Dplus[3737] = 14'b0000000_0000000;
		Dplus[3738] = 14'b0000000_0000000;
		Dplus[3739] = 14'b0000000_0000000;
		Dplus[3740] = 14'b0000000_0000000;
		Dplus[3741] = 14'b0000000_0000000;
		Dplus[3742] = 14'b0000000_0000000;
		Dplus[3743] = 14'b0000000_0000000;
		Dplus[3744] = 14'b0000000_0000000;
		Dplus[3745] = 14'b0000000_0000000;
		Dplus[3746] = 14'b0000000_0000000;
		Dplus[3747] = 14'b0000000_0000000;
		Dplus[3748] = 14'b0000000_0000000;
		Dplus[3749] = 14'b0000000_0000000;
		Dplus[3750] = 14'b0000000_0000000;
		Dplus[3751] = 14'b0000000_0000000;
		Dplus[3752] = 14'b0000000_0000000;
		Dplus[3753] = 14'b0000000_0000000;
		Dplus[3754] = 14'b0000000_0000000;
		Dplus[3755] = 14'b0000000_0000000;
		Dplus[3756] = 14'b0000000_0000000;
		Dplus[3757] = 14'b0000000_0000000;
		Dplus[3758] = 14'b0000000_0000000;
		Dplus[3759] = 14'b0000000_0000000;
		Dplus[3760] = 14'b0000000_0000000;
		Dplus[3761] = 14'b0000000_0000000;
		Dplus[3762] = 14'b0000000_0000000;
		Dplus[3763] = 14'b0000000_0000000;
		Dplus[3764] = 14'b0000000_0000000;
		Dplus[3765] = 14'b0000000_0000000;
		Dplus[3766] = 14'b0000000_0000000;
		Dplus[3767] = 14'b0000000_0000000;
		Dplus[3768] = 14'b0000000_0000000;
		Dplus[3769] = 14'b0000000_0000000;
		Dplus[3770] = 14'b0000000_0000000;
		Dplus[3771] = 14'b0000000_0000000;
		Dplus[3772] = 14'b0000000_0000000;
		Dplus[3773] = 14'b0000000_0000000;
		Dplus[3774] = 14'b0000000_0000000;
		Dplus[3775] = 14'b0000000_0000000;
		Dplus[3776] = 14'b0000000_0000000;
		Dplus[3777] = 14'b0000000_0000000;
		Dplus[3778] = 14'b0000000_0000000;
		Dplus[3779] = 14'b0000000_0000000;
		Dplus[3780] = 14'b0000000_0000000;
		Dplus[3781] = 14'b0000000_0000000;
		Dplus[3782] = 14'b0000000_0000000;
		Dplus[3783] = 14'b0000000_0000000;
		Dplus[3784] = 14'b0000000_0000000;
		Dplus[3785] = 14'b0000000_0000000;
		Dplus[3786] = 14'b0000000_0000000;
		Dplus[3787] = 14'b0000000_0000000;
		Dplus[3788] = 14'b0000000_0000000;
		Dplus[3789] = 14'b0000000_0000000;
		Dplus[3790] = 14'b0000000_0000000;
		Dplus[3791] = 14'b0000000_0000000;
		Dplus[3792] = 14'b0000000_0000000;
		Dplus[3793] = 14'b0000000_0000000;
		Dplus[3794] = 14'b0000000_0000000;
		Dplus[3795] = 14'b0000000_0000000;
		Dplus[3796] = 14'b0000000_0000000;
		Dplus[3797] = 14'b0000000_0000000;
		Dplus[3798] = 14'b0000000_0000000;
		Dplus[3799] = 14'b0000000_0000000;
		Dplus[3800] = 14'b0000000_0000000;
		Dplus[3801] = 14'b0000000_0000000;
		Dplus[3802] = 14'b0000000_0000000;
		Dplus[3803] = 14'b0000000_0000000;
		Dplus[3804] = 14'b0000000_0000000;
		Dplus[3805] = 14'b0000000_0000000;
		Dplus[3806] = 14'b0000000_0000000;
		Dplus[3807] = 14'b0000000_0000000;
		Dplus[3808] = 14'b0000000_0000000;
		Dplus[3809] = 14'b0000000_0000000;
		Dplus[3810] = 14'b0000000_0000000;
		Dplus[3811] = 14'b0000000_0000000;
		Dplus[3812] = 14'b0000000_0000000;
		Dplus[3813] = 14'b0000000_0000000;
		Dplus[3814] = 14'b0000000_0000000;
		Dplus[3815] = 14'b0000000_0000000;
		Dplus[3816] = 14'b0000000_0000000;
		Dplus[3817] = 14'b0000000_0000000;
		Dplus[3818] = 14'b0000000_0000000;
		Dplus[3819] = 14'b0000000_0000000;
		Dplus[3820] = 14'b0000000_0000000;
		Dplus[3821] = 14'b0000000_0000000;
		Dplus[3822] = 14'b0000000_0000000;
		Dplus[3823] = 14'b0000000_0000000;
		Dplus[3824] = 14'b0000000_0000000;
		Dplus[3825] = 14'b0000000_0000000;
		Dplus[3826] = 14'b0000000_0000000;
		Dplus[3827] = 14'b0000000_0000000;
		Dplus[3828] = 14'b0000000_0000000;
		Dplus[3829] = 14'b0000000_0000000;
		Dplus[3830] = 14'b0000000_0000000;
		Dplus[3831] = 14'b0000000_0000000;
		Dplus[3832] = 14'b0000000_0000000;
		Dplus[3833] = 14'b0000000_0000000;
		Dplus[3834] = 14'b0000000_0000000;
		Dplus[3835] = 14'b0000000_0000000;
		Dplus[3836] = 14'b0000000_0000000;
		Dplus[3837] = 14'b0000000_0000000;
		Dplus[3838] = 14'b0000000_0000000;
		Dplus[3839] = 14'b0000000_0000000;
		Dplus[3840] = 14'b0000000_0000000;
		Dplus[3841] = 14'b0000000_0000000;
		Dplus[3842] = 14'b0000000_0000000;
		Dplus[3843] = 14'b0000000_0000000;
		Dplus[3844] = 14'b0000000_0000000;
		Dplus[3845] = 14'b0000000_0000000;
		Dplus[3846] = 14'b0000000_0000000;
		Dplus[3847] = 14'b0000000_0000000;
		Dplus[3848] = 14'b0000000_0000000;
		Dplus[3849] = 14'b0000000_0000000;
		Dplus[3850] = 14'b0000000_0000000;
		Dplus[3851] = 14'b0000000_0000000;
		Dplus[3852] = 14'b0000000_0000000;
		Dplus[3853] = 14'b0000000_0000000;
		Dplus[3854] = 14'b0000000_0000000;
		Dplus[3855] = 14'b0000000_0000000;
		Dplus[3856] = 14'b0000000_0000000;
		Dplus[3857] = 14'b0000000_0000000;
		Dplus[3858] = 14'b0000000_0000000;
		Dplus[3859] = 14'b0000000_0000000;
		Dplus[3860] = 14'b0000000_0000000;
		Dplus[3861] = 14'b0000000_0000000;
		Dplus[3862] = 14'b0000000_0000000;
		Dplus[3863] = 14'b0000000_0000000;
		Dplus[3864] = 14'b0000000_0000000;
		Dplus[3865] = 14'b0000000_0000000;
		Dplus[3866] = 14'b0000000_0000000;
		Dplus[3867] = 14'b0000000_0000000;
		Dplus[3868] = 14'b0000000_0000000;
		Dplus[3869] = 14'b0000000_0000000;
		Dplus[3870] = 14'b0000000_0000000;
		Dplus[3871] = 14'b0000000_0000000;
		Dplus[3872] = 14'b0000000_0000000;
		Dplus[3873] = 14'b0000000_0000000;
		Dplus[3874] = 14'b0000000_0000000;
		Dplus[3875] = 14'b0000000_0000000;
		Dplus[3876] = 14'b0000000_0000000;
		Dplus[3877] = 14'b0000000_0000000;
		Dplus[3878] = 14'b0000000_0000000;
		Dplus[3879] = 14'b0000000_0000000;
		Dplus[3880] = 14'b0000000_0000000;
		Dplus[3881] = 14'b0000000_0000000;
		Dplus[3882] = 14'b0000000_0000000;
		Dplus[3883] = 14'b0000000_0000000;
		Dplus[3884] = 14'b0000000_0000000;
		Dplus[3885] = 14'b0000000_0000000;
		Dplus[3886] = 14'b0000000_0000000;
		Dplus[3887] = 14'b0000000_0000000;
		Dplus[3888] = 14'b0000000_0000000;
		Dplus[3889] = 14'b0000000_0000000;
		Dplus[3890] = 14'b0000000_0000000;
		Dplus[3891] = 14'b0000000_0000000;
		Dplus[3892] = 14'b0000000_0000000;
		Dplus[3893] = 14'b0000000_0000000;
		Dplus[3894] = 14'b0000000_0000000;
		Dplus[3895] = 14'b0000000_0000000;
		Dplus[3896] = 14'b0000000_0000000;
		Dplus[3897] = 14'b0000000_0000000;
		Dplus[3898] = 14'b0000000_0000000;
		Dplus[3899] = 14'b0000000_0000000;
		Dplus[3900] = 14'b0000000_0000000;
		Dplus[3901] = 14'b0000000_0000000;
		Dplus[3902] = 14'b0000000_0000000;
		Dplus[3903] = 14'b0000000_0000000;
		Dplus[3904] = 14'b0000000_0000000;
		Dplus[3905] = 14'b0000000_0000000;
		Dplus[3906] = 14'b0000000_0000000;
		Dplus[3907] = 14'b0000000_0000000;
		Dplus[3908] = 14'b0000000_0000000;
		Dplus[3909] = 14'b0000000_0000000;
		Dplus[3910] = 14'b0000000_0000000;
		Dplus[3911] = 14'b0000000_0000000;
		Dplus[3912] = 14'b0000000_0000000;
		Dplus[3913] = 14'b0000000_0000000;
		Dplus[3914] = 14'b0000000_0000000;
		Dplus[3915] = 14'b0000000_0000000;
		Dplus[3916] = 14'b0000000_0000000;
		Dplus[3917] = 14'b0000000_0000000;
		Dplus[3918] = 14'b0000000_0000000;
		Dplus[3919] = 14'b0000000_0000000;
		Dplus[3920] = 14'b0000000_0000000;
		Dplus[3921] = 14'b0000000_0000000;
		Dplus[3922] = 14'b0000000_0000000;
		Dplus[3923] = 14'b0000000_0000000;
		Dplus[3924] = 14'b0000000_0000000;
		Dplus[3925] = 14'b0000000_0000000;
		Dplus[3926] = 14'b0000000_0000000;
		Dplus[3927] = 14'b0000000_0000000;
		Dplus[3928] = 14'b0000000_0000000;
		Dplus[3929] = 14'b0000000_0000000;
		Dplus[3930] = 14'b0000000_0000000;
		Dplus[3931] = 14'b0000000_0000000;
		Dplus[3932] = 14'b0000000_0000000;
		Dplus[3933] = 14'b0000000_0000000;
		Dplus[3934] = 14'b0000000_0000000;
		Dplus[3935] = 14'b0000000_0000000;
		Dplus[3936] = 14'b0000000_0000000;
		Dplus[3937] = 14'b0000000_0000000;
		Dplus[3938] = 14'b0000000_0000000;
		Dplus[3939] = 14'b0000000_0000000;
		Dplus[3940] = 14'b0000000_0000000;
		Dplus[3941] = 14'b0000000_0000000;
		Dplus[3942] = 14'b0000000_0000000;
		Dplus[3943] = 14'b0000000_0000000;
		Dplus[3944] = 14'b0000000_0000000;
		Dplus[3945] = 14'b0000000_0000000;
		Dplus[3946] = 14'b0000000_0000000;
		Dplus[3947] = 14'b0000000_0000000;
		Dplus[3948] = 14'b0000000_0000000;
		Dplus[3949] = 14'b0000000_0000000;
		Dplus[3950] = 14'b0000000_0000000;
		Dplus[3951] = 14'b0000000_0000000;
		Dplus[3952] = 14'b0000000_0000000;
		Dplus[3953] = 14'b0000000_0000000;
		Dplus[3954] = 14'b0000000_0000000;
		Dplus[3955] = 14'b0000000_0000000;
		Dplus[3956] = 14'b0000000_0000000;
		Dplus[3957] = 14'b0000000_0000000;
		Dplus[3958] = 14'b0000000_0000000;
		Dplus[3959] = 14'b0000000_0000000;
		Dplus[3960] = 14'b0000000_0000000;
		Dplus[3961] = 14'b0000000_0000000;
		Dplus[3962] = 14'b0000000_0000000;
		Dplus[3963] = 14'b0000000_0000000;
		Dplus[3964] = 14'b0000000_0000000;
		Dplus[3965] = 14'b0000000_0000000;
		Dplus[3966] = 14'b0000000_0000000;
		Dplus[3967] = 14'b0000000_0000000;
		Dplus[3968] = 14'b0000000_0000000;
		Dplus[3969] = 14'b0000000_0000000;
		Dplus[3970] = 14'b0000000_0000000;
		Dplus[3971] = 14'b0000000_0000000;
		Dplus[3972] = 14'b0000000_0000000;
		Dplus[3973] = 14'b0000000_0000000;
		Dplus[3974] = 14'b0000000_0000000;
		Dplus[3975] = 14'b0000000_0000000;
		Dplus[3976] = 14'b0000000_0000000;
		Dplus[3977] = 14'b0000000_0000000;
		Dplus[3978] = 14'b0000000_0000000;
		Dplus[3979] = 14'b0000000_0000000;
		Dplus[3980] = 14'b0000000_0000000;
		Dplus[3981] = 14'b0000000_0000000;
		Dplus[3982] = 14'b0000000_0000000;
		Dplus[3983] = 14'b0000000_0000000;
		Dplus[3984] = 14'b0000000_0000000;
		Dplus[3985] = 14'b0000000_0000000;
		Dplus[3986] = 14'b0000000_0000000;
		Dplus[3987] = 14'b0000000_0000000;
		Dplus[3988] = 14'b0000000_0000000;
		Dplus[3989] = 14'b0000000_0000000;
		Dplus[3990] = 14'b0000000_0000000;
		Dplus[3991] = 14'b0000000_0000000;
		Dplus[3992] = 14'b0000000_0000000;
		Dplus[3993] = 14'b0000000_0000000;
		Dplus[3994] = 14'b0000000_0000000;
		Dplus[3995] = 14'b0000000_0000000;
		Dplus[3996] = 14'b0000000_0000000;
		Dplus[3997] = 14'b0000000_0000000;
		Dplus[3998] = 14'b0000000_0000000;
		Dplus[3999] = 14'b0000000_0000000;
		Dplus[4000] = 14'b0000000_0000000;
		Dplus[4001] = 14'b0000000_0000000;
		Dplus[4002] = 14'b0000000_0000000;
		Dplus[4003] = 14'b0000000_0000000;
		Dplus[4004] = 14'b0000000_0000000;
		Dplus[4005] = 14'b0000000_0000000;
		Dplus[4006] = 14'b0000000_0000000;
		Dplus[4007] = 14'b0000000_0000000;
		Dplus[4008] = 14'b0000000_0000000;
		Dplus[4009] = 14'b0000000_0000000;
		Dplus[4010] = 14'b0000000_0000000;
		Dplus[4011] = 14'b0000000_0000000;
		Dplus[4012] = 14'b0000000_0000000;
		Dplus[4013] = 14'b0000000_0000000;
		Dplus[4014] = 14'b0000000_0000000;
		Dplus[4015] = 14'b0000000_0000000;
		Dplus[4016] = 14'b0000000_0000000;
		Dplus[4017] = 14'b0000000_0000000;
		Dplus[4018] = 14'b0000000_0000000;
		Dplus[4019] = 14'b0000000_0000000;
		Dplus[4020] = 14'b0000000_0000000;
		Dplus[4021] = 14'b0000000_0000000;
		Dplus[4022] = 14'b0000000_0000000;
		Dplus[4023] = 14'b0000000_0000000;
		Dplus[4024] = 14'b0000000_0000000;
		Dplus[4025] = 14'b0000000_0000000;
		Dplus[4026] = 14'b0000000_0000000;
		Dplus[4027] = 14'b0000000_0000000;
		Dplus[4028] = 14'b0000000_0000000;
		Dplus[4029] = 14'b0000000_0000000;
		Dplus[4030] = 14'b0000000_0000000;
		Dplus[4031] = 14'b0000000_0000000;
		Dplus[4032] = 14'b0000000_0000000;
		Dplus[4033] = 14'b0000000_0000000;
		Dplus[4034] = 14'b0000000_0000000;
		Dplus[4035] = 14'b0000000_0000000;
		Dplus[4036] = 14'b0000000_0000000;
		Dplus[4037] = 14'b0000000_0000000;
		Dplus[4038] = 14'b0000000_0000000;
		Dplus[4039] = 14'b0000000_0000000;
		Dplus[4040] = 14'b0000000_0000000;
		Dplus[4041] = 14'b0000000_0000000;
		Dplus[4042] = 14'b0000000_0000000;
		Dplus[4043] = 14'b0000000_0000000;
		Dplus[4044] = 14'b0000000_0000000;
		Dplus[4045] = 14'b0000000_0000000;
		Dplus[4046] = 14'b0000000_0000000;
		Dplus[4047] = 14'b0000000_0000000;
		Dplus[4048] = 14'b0000000_0000000;
		Dplus[4049] = 14'b0000000_0000000;
		Dplus[4050] = 14'b0000000_0000000;
		Dplus[4051] = 14'b0000000_0000000;
		Dplus[4052] = 14'b0000000_0000000;
		Dplus[4053] = 14'b0000000_0000000;
		Dplus[4054] = 14'b0000000_0000000;
		Dplus[4055] = 14'b0000000_0000000;
		Dplus[4056] = 14'b0000000_0000000;
		Dplus[4057] = 14'b0000000_0000000;
		Dplus[4058] = 14'b0000000_0000000;
		Dplus[4059] = 14'b0000000_0000000;
		Dplus[4060] = 14'b0000000_0000000;
		Dplus[4061] = 14'b0000000_0000000;
		Dplus[4062] = 14'b0000000_0000000;
		Dplus[4063] = 14'b0000000_0000000;
		Dplus[4064] = 14'b0000000_0000000;
		Dplus[4065] = 14'b0000000_0000000;
		Dplus[4066] = 14'b0000000_0000000;
		Dplus[4067] = 14'b0000000_0000000;
		Dplus[4068] = 14'b0000000_0000000;
		Dplus[4069] = 14'b0000000_0000000;
		Dplus[4070] = 14'b0000000_0000000;
		Dplus[4071] = 14'b0000000_0000000;
		Dplus[4072] = 14'b0000000_0000000;
		Dplus[4073] = 14'b0000000_0000000;
		Dplus[4074] = 14'b0000000_0000000;
		Dplus[4075] = 14'b0000000_0000000;
		Dplus[4076] = 14'b0000000_0000000;
		Dplus[4077] = 14'b0000000_0000000;
		Dplus[4078] = 14'b0000000_0000000;
		Dplus[4079] = 14'b0000000_0000000;
		Dplus[4080] = 14'b0000000_0000000;
		Dplus[4081] = 14'b0000000_0000000;
		Dplus[4082] = 14'b0000000_0000000;
		Dplus[4083] = 14'b0000000_0000000;
		Dplus[4084] = 14'b0000000_0000000;
		Dplus[4085] = 14'b0000000_0000000;
		Dplus[4086] = 14'b0000000_0000000;
		Dplus[4087] = 14'b0000000_0000000;
		Dplus[4088] = 14'b0000000_0000000;
		Dplus[4089] = 14'b0000000_0000000;
		Dplus[4090] = 14'b0000000_0000000;
		Dplus[4091] = 14'b0000000_0000000;
		Dplus[4092] = 14'b0000000_0000000;
		Dplus[4093] = 14'b0000000_0000000;
		Dplus[4094] = 14'b0000000_0000000;
		Dplus[4095] = 14'b0000000_0000000;
		Dplus[4096] = 14'b0000000_0000000;
		Dplus[4097] = 14'b0000000_0000000;
		Dplus[4098] = 14'b0000000_0000000;
		Dplus[4099] = 14'b0000000_0000000;
		Dplus[4100] = 14'b0000000_0000000;
		Dplus[4101] = 14'b0000000_0000000;
		Dplus[4102] = 14'b0000000_0000000;
		Dplus[4103] = 14'b0000000_0000000;
		Dplus[4104] = 14'b0000000_0000000;
		Dplus[4105] = 14'b0000000_0000000;
		Dplus[4106] = 14'b0000000_0000000;
		Dplus[4107] = 14'b0000000_0000000;
		Dplus[4108] = 14'b0000000_0000000;
		Dplus[4109] = 14'b0000000_0000000;
		Dplus[4110] = 14'b0000000_0000000;
		Dplus[4111] = 14'b0000000_0000000;
		Dplus[4112] = 14'b0000000_0000000;
		Dplus[4113] = 14'b0000000_0000000;
		Dplus[4114] = 14'b0000000_0000000;
		Dplus[4115] = 14'b0000000_0000000;
		Dplus[4116] = 14'b0000000_0000000;
		Dplus[4117] = 14'b0000000_0000000;
		Dplus[4118] = 14'b0000000_0000000;
		Dplus[4119] = 14'b0000000_0000000;
		Dplus[4120] = 14'b0000000_0000000;
		Dplus[4121] = 14'b0000000_0000000;
		Dplus[4122] = 14'b0000000_0000000;
		Dplus[4123] = 14'b0000000_0000000;
		Dplus[4124] = 14'b0000000_0000000;
		Dplus[4125] = 14'b0000000_0000000;
		Dplus[4126] = 14'b0000000_0000000;
		Dplus[4127] = 14'b0000000_0000000;
		Dplus[4128] = 14'b0000000_0000000;
		Dplus[4129] = 14'b0000000_0000000;
		Dplus[4130] = 14'b0000000_0000000;
		Dplus[4131] = 14'b0000000_0000000;
		Dplus[4132] = 14'b0000000_0000000;
		Dplus[4133] = 14'b0000000_0000000;
		Dplus[4134] = 14'b0000000_0000000;
		Dplus[4135] = 14'b0000000_0000000;
		Dplus[4136] = 14'b0000000_0000000;
		Dplus[4137] = 14'b0000000_0000000;
		Dplus[4138] = 14'b0000000_0000000;
		Dplus[4139] = 14'b0000000_0000000;
		Dplus[4140] = 14'b0000000_0000000;
		Dplus[4141] = 14'b0000000_0000000;
		Dplus[4142] = 14'b0000000_0000000;
		Dplus[4143] = 14'b0000000_0000000;
		Dplus[4144] = 14'b0000000_0000000;
		Dplus[4145] = 14'b0000000_0000000;
		Dplus[4146] = 14'b0000000_0000000;
		Dplus[4147] = 14'b0000000_0000000;
		Dplus[4148] = 14'b0000000_0000000;
		Dplus[4149] = 14'b0000000_0000000;
		Dplus[4150] = 14'b0000000_0000000;
		Dplus[4151] = 14'b0000000_0000000;
		Dplus[4152] = 14'b0000000_0000000;
		Dplus[4153] = 14'b0000000_0000000;
		Dplus[4154] = 14'b0000000_0000000;
		Dplus[4155] = 14'b0000000_0000000;
		Dplus[4156] = 14'b0000000_0000000;
		Dplus[4157] = 14'b0000000_0000000;
		Dplus[4158] = 14'b0000000_0000000;
		Dplus[4159] = 14'b0000000_0000000;
		Dplus[4160] = 14'b0000000_0000000;
		Dplus[4161] = 14'b0000000_0000000;
		Dplus[4162] = 14'b0000000_0000000;
		Dplus[4163] = 14'b0000000_0000000;
		Dplus[4164] = 14'b0000000_0000000;
		Dplus[4165] = 14'b0000000_0000000;
		Dplus[4166] = 14'b0000000_0000000;
		Dplus[4167] = 14'b0000000_0000000;
		Dplus[4168] = 14'b0000000_0000000;
		Dplus[4169] = 14'b0000000_0000000;
		Dplus[4170] = 14'b0000000_0000000;
		Dplus[4171] = 14'b0000000_0000000;
		Dplus[4172] = 14'b0000000_0000000;
		Dplus[4173] = 14'b0000000_0000000;
		Dplus[4174] = 14'b0000000_0000000;
		Dplus[4175] = 14'b0000000_0000000;
		Dplus[4176] = 14'b0000000_0000000;
		Dplus[4177] = 14'b0000000_0000000;
		Dplus[4178] = 14'b0000000_0000000;
		Dplus[4179] = 14'b0000000_0000000;
		Dplus[4180] = 14'b0000000_0000000;
		Dplus[4181] = 14'b0000000_0000000;
		Dplus[4182] = 14'b0000000_0000000;
		Dplus[4183] = 14'b0000000_0000000;
		Dplus[4184] = 14'b0000000_0000000;
		Dplus[4185] = 14'b0000000_0000000;
		Dplus[4186] = 14'b0000000_0000000;
		Dplus[4187] = 14'b0000000_0000000;
		Dplus[4188] = 14'b0000000_0000000;
		Dplus[4189] = 14'b0000000_0000000;
		Dplus[4190] = 14'b0000000_0000000;
		Dplus[4191] = 14'b0000000_0000000;
		Dplus[4192] = 14'b0000000_0000000;
		Dplus[4193] = 14'b0000000_0000000;
		Dplus[4194] = 14'b0000000_0000000;
		Dplus[4195] = 14'b0000000_0000000;
		Dplus[4196] = 14'b0000000_0000000;
		Dplus[4197] = 14'b0000000_0000000;
		Dplus[4198] = 14'b0000000_0000000;
		Dplus[4199] = 14'b0000000_0000000;
		Dplus[4200] = 14'b0000000_0000000;
		Dplus[4201] = 14'b0000000_0000000;
		Dplus[4202] = 14'b0000000_0000000;
		Dplus[4203] = 14'b0000000_0000000;
		Dplus[4204] = 14'b0000000_0000000;
		Dplus[4205] = 14'b0000000_0000000;
		Dplus[4206] = 14'b0000000_0000000;
		Dplus[4207] = 14'b0000000_0000000;
		Dplus[4208] = 14'b0000000_0000000;
		Dplus[4209] = 14'b0000000_0000000;
		Dplus[4210] = 14'b0000000_0000000;
		Dplus[4211] = 14'b0000000_0000000;
		Dplus[4212] = 14'b0000000_0000000;
		Dplus[4213] = 14'b0000000_0000000;
		Dplus[4214] = 14'b0000000_0000000;
		Dplus[4215] = 14'b0000000_0000000;
		Dplus[4216] = 14'b0000000_0000000;
		Dplus[4217] = 14'b0000000_0000000;
		Dplus[4218] = 14'b0000000_0000000;
		Dplus[4219] = 14'b0000000_0000000;
		Dplus[4220] = 14'b0000000_0000000;
		Dplus[4221] = 14'b0000000_0000000;
		Dplus[4222] = 14'b0000000_0000000;
		Dplus[4223] = 14'b0000000_0000000;
		Dplus[4224] = 14'b0000000_0000000;
		Dplus[4225] = 14'b0000000_0000000;
		Dplus[4226] = 14'b0000000_0000000;
		Dplus[4227] = 14'b0000000_0000000;
		Dplus[4228] = 14'b0000000_0000000;
		Dplus[4229] = 14'b0000000_0000000;
		Dplus[4230] = 14'b0000000_0000000;
		Dplus[4231] = 14'b0000000_0000000;
		Dplus[4232] = 14'b0000000_0000000;
		Dplus[4233] = 14'b0000000_0000000;
		Dplus[4234] = 14'b0000000_0000000;
		Dplus[4235] = 14'b0000000_0000000;
		Dplus[4236] = 14'b0000000_0000000;
		Dplus[4237] = 14'b0000000_0000000;
		Dplus[4238] = 14'b0000000_0000000;
		Dplus[4239] = 14'b0000000_0000000;
		Dplus[4240] = 14'b0000000_0000000;
		Dplus[4241] = 14'b0000000_0000000;
		Dplus[4242] = 14'b0000000_0000000;
		Dplus[4243] = 14'b0000000_0000000;
		Dplus[4244] = 14'b0000000_0000000;
		Dplus[4245] = 14'b0000000_0000000;
		Dplus[4246] = 14'b0000000_0000000;
		Dplus[4247] = 14'b0000000_0000000;
		Dplus[4248] = 14'b0000000_0000000;
		Dplus[4249] = 14'b0000000_0000000;
		Dplus[4250] = 14'b0000000_0000000;
		Dplus[4251] = 14'b0000000_0000000;
		Dplus[4252] = 14'b0000000_0000000;
		Dplus[4253] = 14'b0000000_0000000;
		Dplus[4254] = 14'b0000000_0000000;
		Dplus[4255] = 14'b0000000_0000000;
		Dplus[4256] = 14'b0000000_0000000;
		Dplus[4257] = 14'b0000000_0000000;
		Dplus[4258] = 14'b0000000_0000000;
		Dplus[4259] = 14'b0000000_0000000;
		Dplus[4260] = 14'b0000000_0000000;
		Dplus[4261] = 14'b0000000_0000000;
		Dplus[4262] = 14'b0000000_0000000;
		Dplus[4263] = 14'b0000000_0000000;
		Dplus[4264] = 14'b0000000_0000000;
		Dplus[4265] = 14'b0000000_0000000;
		Dplus[4266] = 14'b0000000_0000000;
		Dplus[4267] = 14'b0000000_0000000;
		Dplus[4268] = 14'b0000000_0000000;
		Dplus[4269] = 14'b0000000_0000000;
		Dplus[4270] = 14'b0000000_0000000;
		Dplus[4271] = 14'b0000000_0000000;
		Dplus[4272] = 14'b0000000_0000000;
		Dplus[4273] = 14'b0000000_0000000;
		Dplus[4274] = 14'b0000000_0000000;
		Dplus[4275] = 14'b0000000_0000000;
		Dplus[4276] = 14'b0000000_0000000;
		Dplus[4277] = 14'b0000000_0000000;
		Dplus[4278] = 14'b0000000_0000000;
		Dplus[4279] = 14'b0000000_0000000;
		Dplus[4280] = 14'b0000000_0000000;
		Dplus[4281] = 14'b0000000_0000000;
		Dplus[4282] = 14'b0000000_0000000;
		Dplus[4283] = 14'b0000000_0000000;
		Dplus[4284] = 14'b0000000_0000000;
		Dplus[4285] = 14'b0000000_0000000;
		Dplus[4286] = 14'b0000000_0000000;
		Dplus[4287] = 14'b0000000_0000000;
		Dplus[4288] = 14'b0000000_0000000;
		Dplus[4289] = 14'b0000000_0000000;
		Dplus[4290] = 14'b0000000_0000000;
		Dplus[4291] = 14'b0000000_0000000;
		Dplus[4292] = 14'b0000000_0000000;
		Dplus[4293] = 14'b0000000_0000000;
		Dplus[4294] = 14'b0000000_0000000;
		Dplus[4295] = 14'b0000000_0000000;
		Dplus[4296] = 14'b0000000_0000000;
		Dplus[4297] = 14'b0000000_0000000;
		Dplus[4298] = 14'b0000000_0000000;
		Dplus[4299] = 14'b0000000_0000000;
		Dplus[4300] = 14'b0000000_0000000;
		Dplus[4301] = 14'b0000000_0000000;
		Dplus[4302] = 14'b0000000_0000000;
		Dplus[4303] = 14'b0000000_0000000;
		Dplus[4304] = 14'b0000000_0000000;
		Dplus[4305] = 14'b0000000_0000000;
		Dplus[4306] = 14'b0000000_0000000;
		Dplus[4307] = 14'b0000000_0000000;
		Dplus[4308] = 14'b0000000_0000000;
		Dplus[4309] = 14'b0000000_0000000;
		Dplus[4310] = 14'b0000000_0000000;
		Dplus[4311] = 14'b0000000_0000000;
		Dplus[4312] = 14'b0000000_0000000;
		Dplus[4313] = 14'b0000000_0000000;
		Dplus[4314] = 14'b0000000_0000000;
		Dplus[4315] = 14'b0000000_0000000;
		Dplus[4316] = 14'b0000000_0000000;
		Dplus[4317] = 14'b0000000_0000000;
		Dplus[4318] = 14'b0000000_0000000;
		Dplus[4319] = 14'b0000000_0000000;
		Dplus[4320] = 14'b0000000_0000000;
		Dplus[4321] = 14'b0000000_0000000;
		Dplus[4322] = 14'b0000000_0000000;
		Dplus[4323] = 14'b0000000_0000000;
		Dplus[4324] = 14'b0000000_0000000;
		Dplus[4325] = 14'b0000000_0000000;
		Dplus[4326] = 14'b0000000_0000000;
		Dplus[4327] = 14'b0000000_0000000;
		Dplus[4328] = 14'b0000000_0000000;
		Dplus[4329] = 14'b0000000_0000000;
		Dplus[4330] = 14'b0000000_0000000;
		Dplus[4331] = 14'b0000000_0000000;
		Dplus[4332] = 14'b0000000_0000000;
		Dplus[4333] = 14'b0000000_0000000;
		Dplus[4334] = 14'b0000000_0000000;
		Dplus[4335] = 14'b0000000_0000000;
		Dplus[4336] = 14'b0000000_0000000;
		Dplus[4337] = 14'b0000000_0000000;
		Dplus[4338] = 14'b0000000_0000000;
		Dplus[4339] = 14'b0000000_0000000;
		Dplus[4340] = 14'b0000000_0000000;
		Dplus[4341] = 14'b0000000_0000000;
		Dplus[4342] = 14'b0000000_0000000;
		Dplus[4343] = 14'b0000000_0000000;
		Dplus[4344] = 14'b0000000_0000000;
		Dplus[4345] = 14'b0000000_0000000;
		Dplus[4346] = 14'b0000000_0000000;
		Dplus[4347] = 14'b0000000_0000000;
		Dplus[4348] = 14'b0000000_0000000;
		Dplus[4349] = 14'b0000000_0000000;
		Dplus[4350] = 14'b0000000_0000000;
		Dplus[4351] = 14'b0000000_0000000;
		Dplus[4352] = 14'b0000000_0000000;
		Dplus[4353] = 14'b0000000_0000000;
		Dplus[4354] = 14'b0000000_0000000;
		Dplus[4355] = 14'b0000000_0000000;
		Dplus[4356] = 14'b0000000_0000000;
		Dplus[4357] = 14'b0000000_0000000;
		Dplus[4358] = 14'b0000000_0000000;
		Dplus[4359] = 14'b0000000_0000000;
		Dplus[4360] = 14'b0000000_0000000;
		Dplus[4361] = 14'b0000000_0000000;
		Dplus[4362] = 14'b0000000_0000000;
		Dplus[4363] = 14'b0000000_0000000;
		Dplus[4364] = 14'b0000000_0000000;
		Dplus[4365] = 14'b0000000_0000000;
		Dplus[4366] = 14'b0000000_0000000;
		Dplus[4367] = 14'b0000000_0000000;
		Dplus[4368] = 14'b0000000_0000000;
		Dplus[4369] = 14'b0000000_0000000;
		Dplus[4370] = 14'b0000000_0000000;
		Dplus[4371] = 14'b0000000_0000000;
		Dplus[4372] = 14'b0000000_0000000;
		Dplus[4373] = 14'b0000000_0000000;
		Dplus[4374] = 14'b0000000_0000000;
		Dplus[4375] = 14'b0000000_0000000;
		Dplus[4376] = 14'b0000000_0000000;
		Dplus[4377] = 14'b0000000_0000000;
		Dplus[4378] = 14'b0000000_0000000;
		Dplus[4379] = 14'b0000000_0000000;
		Dplus[4380] = 14'b0000000_0000000;
		Dplus[4381] = 14'b0000000_0000000;
		Dplus[4382] = 14'b0000000_0000000;
		Dplus[4383] = 14'b0000000_0000000;
		Dplus[4384] = 14'b0000000_0000000;
		Dplus[4385] = 14'b0000000_0000000;
		Dplus[4386] = 14'b0000000_0000000;
		Dplus[4387] = 14'b0000000_0000000;
		Dplus[4388] = 14'b0000000_0000000;
		Dplus[4389] = 14'b0000000_0000000;
		Dplus[4390] = 14'b0000000_0000000;
		Dplus[4391] = 14'b0000000_0000000;
		Dplus[4392] = 14'b0000000_0000000;
		Dplus[4393] = 14'b0000000_0000000;
		Dplus[4394] = 14'b0000000_0000000;
		Dplus[4395] = 14'b0000000_0000000;
		Dplus[4396] = 14'b0000000_0000000;
		Dplus[4397] = 14'b0000000_0000000;
		Dplus[4398] = 14'b0000000_0000000;
		Dplus[4399] = 14'b0000000_0000000;
		Dplus[4400] = 14'b0000000_0000000;
		Dplus[4401] = 14'b0000000_0000000;
		Dplus[4402] = 14'b0000000_0000000;
		Dplus[4403] = 14'b0000000_0000000;
		Dplus[4404] = 14'b0000000_0000000;
		Dplus[4405] = 14'b0000000_0000000;
		Dplus[4406] = 14'b0000000_0000000;
		Dplus[4407] = 14'b0000000_0000000;
		Dplus[4408] = 14'b0000000_0000000;
		Dplus[4409] = 14'b0000000_0000000;
		Dplus[4410] = 14'b0000000_0000000;
		Dplus[4411] = 14'b0000000_0000000;
		Dplus[4412] = 14'b0000000_0000000;
		Dplus[4413] = 14'b0000000_0000000;
		Dplus[4414] = 14'b0000000_0000000;
		Dplus[4415] = 14'b0000000_0000000;
		Dplus[4416] = 14'b0000000_0000000;
		Dplus[4417] = 14'b0000000_0000000;
		Dplus[4418] = 14'b0000000_0000000;
		Dplus[4419] = 14'b0000000_0000000;
		Dplus[4420] = 14'b0000000_0000000;
		Dplus[4421] = 14'b0000000_0000000;
		Dplus[4422] = 14'b0000000_0000000;
		Dplus[4423] = 14'b0000000_0000000;
		Dplus[4424] = 14'b0000000_0000000;
		Dplus[4425] = 14'b0000000_0000000;
		Dplus[4426] = 14'b0000000_0000000;
		Dplus[4427] = 14'b0000000_0000000;
		Dplus[4428] = 14'b0000000_0000000;
		Dplus[4429] = 14'b0000000_0000000;
		Dplus[4430] = 14'b0000000_0000000;
		Dplus[4431] = 14'b0000000_0000000;
		Dplus[4432] = 14'b0000000_0000000;
		Dplus[4433] = 14'b0000000_0000000;
		Dplus[4434] = 14'b0000000_0000000;
		Dplus[4435] = 14'b0000000_0000000;
		Dplus[4436] = 14'b0000000_0000000;
		Dplus[4437] = 14'b0000000_0000000;
		Dplus[4438] = 14'b0000000_0000000;
		Dplus[4439] = 14'b0000000_0000000;
		Dplus[4440] = 14'b0000000_0000000;
		Dplus[4441] = 14'b0000000_0000000;
		Dplus[4442] = 14'b0000000_0000000;
		Dplus[4443] = 14'b0000000_0000000;
		Dplus[4444] = 14'b0000000_0000000;
		Dplus[4445] = 14'b0000000_0000000;
		Dplus[4446] = 14'b0000000_0000000;
		Dplus[4447] = 14'b0000000_0000000;
		Dplus[4448] = 14'b0000000_0000000;
		Dplus[4449] = 14'b0000000_0000000;
		Dplus[4450] = 14'b0000000_0000000;
		Dplus[4451] = 14'b0000000_0000000;
		Dplus[4452] = 14'b0000000_0000000;
		Dplus[4453] = 14'b0000000_0000000;
		Dplus[4454] = 14'b0000000_0000000;
		Dplus[4455] = 14'b0000000_0000000;
		Dplus[4456] = 14'b0000000_0000000;
		Dplus[4457] = 14'b0000000_0000000;
		Dplus[4458] = 14'b0000000_0000000;
		Dplus[4459] = 14'b0000000_0000000;
		Dplus[4460] = 14'b0000000_0000000;
		Dplus[4461] = 14'b0000000_0000000;
		Dplus[4462] = 14'b0000000_0000000;
		Dplus[4463] = 14'b0000000_0000000;
		Dplus[4464] = 14'b0000000_0000000;
		Dplus[4465] = 14'b0000000_0000000;
		Dplus[4466] = 14'b0000000_0000000;
		Dplus[4467] = 14'b0000000_0000000;
		Dplus[4468] = 14'b0000000_0000000;
		Dplus[4469] = 14'b0000000_0000000;
		Dplus[4470] = 14'b0000000_0000000;
		Dplus[4471] = 14'b0000000_0000000;
		Dplus[4472] = 14'b0000000_0000000;
		Dplus[4473] = 14'b0000000_0000000;
		Dplus[4474] = 14'b0000000_0000000;
		Dplus[4475] = 14'b0000000_0000000;
		Dplus[4476] = 14'b0000000_0000000;
		Dplus[4477] = 14'b0000000_0000000;
		Dplus[4478] = 14'b0000000_0000000;
		Dplus[4479] = 14'b0000000_0000000;
		Dplus[4480] = 14'b0000000_0000000;
		Dplus[4481] = 14'b0000000_0000000;
		Dplus[4482] = 14'b0000000_0000000;
		Dplus[4483] = 14'b0000000_0000000;
		Dplus[4484] = 14'b0000000_0000000;
		Dplus[4485] = 14'b0000000_0000000;
		Dplus[4486] = 14'b0000000_0000000;
		Dplus[4487] = 14'b0000000_0000000;
		Dplus[4488] = 14'b0000000_0000000;
		Dplus[4489] = 14'b0000000_0000000;
		Dplus[4490] = 14'b0000000_0000000;
		Dplus[4491] = 14'b0000000_0000000;
		Dplus[4492] = 14'b0000000_0000000;
		Dplus[4493] = 14'b0000000_0000000;
		Dplus[4494] = 14'b0000000_0000000;
		Dplus[4495] = 14'b0000000_0000000;
		Dplus[4496] = 14'b0000000_0000000;
		Dplus[4497] = 14'b0000000_0000000;
		Dplus[4498] = 14'b0000000_0000000;
		Dplus[4499] = 14'b0000000_0000000;
		Dplus[4500] = 14'b0000000_0000000;
		Dplus[4501] = 14'b0000000_0000000;
		Dplus[4502] = 14'b0000000_0000000;
		Dplus[4503] = 14'b0000000_0000000;
		Dplus[4504] = 14'b0000000_0000000;
		Dplus[4505] = 14'b0000000_0000000;
		Dplus[4506] = 14'b0000000_0000000;
		Dplus[4507] = 14'b0000000_0000000;
		Dplus[4508] = 14'b0000000_0000000;
		Dplus[4509] = 14'b0000000_0000000;
		Dplus[4510] = 14'b0000000_0000000;
		Dplus[4511] = 14'b0000000_0000000;
		Dplus[4512] = 14'b0000000_0000000;
		Dplus[4513] = 14'b0000000_0000000;
		Dplus[4514] = 14'b0000000_0000000;
		Dplus[4515] = 14'b0000000_0000000;
		Dplus[4516] = 14'b0000000_0000000;
		Dplus[4517] = 14'b0000000_0000000;
		Dplus[4518] = 14'b0000000_0000000;
		Dplus[4519] = 14'b0000000_0000000;
		Dplus[4520] = 14'b0000000_0000000;
		Dplus[4521] = 14'b0000000_0000000;
		Dplus[4522] = 14'b0000000_0000000;
		Dplus[4523] = 14'b0000000_0000000;
		Dplus[4524] = 14'b0000000_0000000;
		Dplus[4525] = 14'b0000000_0000000;
		Dplus[4526] = 14'b0000000_0000000;
		Dplus[4527] = 14'b0000000_0000000;
		Dplus[4528] = 14'b0000000_0000000;
		Dplus[4529] = 14'b0000000_0000000;
		Dplus[4530] = 14'b0000000_0000000;
		Dplus[4531] = 14'b0000000_0000000;
		Dplus[4532] = 14'b0000000_0000000;
		Dplus[4533] = 14'b0000000_0000000;
		Dplus[4534] = 14'b0000000_0000000;
		Dplus[4535] = 14'b0000000_0000000;
		Dplus[4536] = 14'b0000000_0000000;
		Dplus[4537] = 14'b0000000_0000000;
		Dplus[4538] = 14'b0000000_0000000;
		Dplus[4539] = 14'b0000000_0000000;
		Dplus[4540] = 14'b0000000_0000000;
		Dplus[4541] = 14'b0000000_0000000;
		Dplus[4542] = 14'b0000000_0000000;
		Dplus[4543] = 14'b0000000_0000000;
		Dplus[4544] = 14'b0000000_0000000;
		Dplus[4545] = 14'b0000000_0000000;
		Dplus[4546] = 14'b0000000_0000000;
		Dplus[4547] = 14'b0000000_0000000;
		Dplus[4548] = 14'b0000000_0000000;
		Dplus[4549] = 14'b0000000_0000000;
		Dplus[4550] = 14'b0000000_0000000;
		Dplus[4551] = 14'b0000000_0000000;
		Dplus[4552] = 14'b0000000_0000000;
		Dplus[4553] = 14'b0000000_0000000;
		Dplus[4554] = 14'b0000000_0000000;
		Dplus[4555] = 14'b0000000_0000000;
		Dplus[4556] = 14'b0000000_0000000;
		Dplus[4557] = 14'b0000000_0000000;
		Dplus[4558] = 14'b0000000_0000000;
		Dplus[4559] = 14'b0000000_0000000;
		Dplus[4560] = 14'b0000000_0000000;
		Dplus[4561] = 14'b0000000_0000000;
		Dplus[4562] = 14'b0000000_0000000;
		Dplus[4563] = 14'b0000000_0000000;
		Dplus[4564] = 14'b0000000_0000000;
		Dplus[4565] = 14'b0000000_0000000;
		Dplus[4566] = 14'b0000000_0000000;
		Dplus[4567] = 14'b0000000_0000000;
		Dplus[4568] = 14'b0000000_0000000;
		Dplus[4569] = 14'b0000000_0000000;
		Dplus[4570] = 14'b0000000_0000000;
		Dplus[4571] = 14'b0000000_0000000;
		Dplus[4572] = 14'b0000000_0000000;
		Dplus[4573] = 14'b0000000_0000000;
		Dplus[4574] = 14'b0000000_0000000;
		Dplus[4575] = 14'b0000000_0000000;
		Dplus[4576] = 14'b0000000_0000000;
		Dplus[4577] = 14'b0000000_0000000;
		Dplus[4578] = 14'b0000000_0000000;
		Dplus[4579] = 14'b0000000_0000000;
		Dplus[4580] = 14'b0000000_0000000;
		Dplus[4581] = 14'b0000000_0000000;
		Dplus[4582] = 14'b0000000_0000000;
		Dplus[4583] = 14'b0000000_0000000;
		Dplus[4584] = 14'b0000000_0000000;
		Dplus[4585] = 14'b0000000_0000000;
		Dplus[4586] = 14'b0000000_0000000;
		Dplus[4587] = 14'b0000000_0000000;
		Dplus[4588] = 14'b0000000_0000000;
		Dplus[4589] = 14'b0000000_0000000;
		Dplus[4590] = 14'b0000000_0000000;
		Dplus[4591] = 14'b0000000_0000000;
		Dplus[4592] = 14'b0000000_0000000;
		Dplus[4593] = 14'b0000000_0000000;
		Dplus[4594] = 14'b0000000_0000000;
		Dplus[4595] = 14'b0000000_0000000;
		Dplus[4596] = 14'b0000000_0000000;
		Dplus[4597] = 14'b0000000_0000000;
		Dplus[4598] = 14'b0000000_0000000;
		Dplus[4599] = 14'b0000000_0000000;
		Dplus[4600] = 14'b0000000_0000000;
		Dplus[4601] = 14'b0000000_0000000;
		Dplus[4602] = 14'b0000000_0000000;
		Dplus[4603] = 14'b0000000_0000000;
		Dplus[4604] = 14'b0000000_0000000;
		Dplus[4605] = 14'b0000000_0000000;
		Dplus[4606] = 14'b0000000_0000000;
		Dplus[4607] = 14'b0000000_0000000;
		Dplus[4608] = 14'b0000000_0000000;
		Dplus[4609] = 14'b0000000_0000000;
		Dplus[4610] = 14'b0000000_0000000;
		Dplus[4611] = 14'b0000000_0000000;
		Dplus[4612] = 14'b0000000_0000000;
		Dplus[4613] = 14'b0000000_0000000;
		Dplus[4614] = 14'b0000000_0000000;
		Dplus[4615] = 14'b0000000_0000000;
		Dplus[4616] = 14'b0000000_0000000;
		Dplus[4617] = 14'b0000000_0000000;
		Dplus[4618] = 14'b0000000_0000000;
		Dplus[4619] = 14'b0000000_0000000;
		Dplus[4620] = 14'b0000000_0000000;
		Dplus[4621] = 14'b0000000_0000000;
		Dplus[4622] = 14'b0000000_0000000;
		Dplus[4623] = 14'b0000000_0000000;
		Dplus[4624] = 14'b0000000_0000000;
		Dplus[4625] = 14'b0000000_0000000;
		Dplus[4626] = 14'b0000000_0000000;
		Dplus[4627] = 14'b0000000_0000000;
		Dplus[4628] = 14'b0000000_0000000;
		Dplus[4629] = 14'b0000000_0000000;
		Dplus[4630] = 14'b0000000_0000000;
		Dplus[4631] = 14'b0000000_0000000;
		Dplus[4632] = 14'b0000000_0000000;
		Dplus[4633] = 14'b0000000_0000000;
		Dplus[4634] = 14'b0000000_0000000;
		Dplus[4635] = 14'b0000000_0000000;
		Dplus[4636] = 14'b0000000_0000000;
		Dplus[4637] = 14'b0000000_0000000;
		Dplus[4638] = 14'b0000000_0000000;
		Dplus[4639] = 14'b0000000_0000000;
		Dplus[4640] = 14'b0000000_0000000;
		Dplus[4641] = 14'b0000000_0000000;
		Dplus[4642] = 14'b0000000_0000000;
		Dplus[4643] = 14'b0000000_0000000;
		Dplus[4644] = 14'b0000000_0000000;
		Dplus[4645] = 14'b0000000_0000000;
		Dplus[4646] = 14'b0000000_0000000;
		Dplus[4647] = 14'b0000000_0000000;
		Dplus[4648] = 14'b0000000_0000000;
		Dplus[4649] = 14'b0000000_0000000;
		Dplus[4650] = 14'b0000000_0000000;
		Dplus[4651] = 14'b0000000_0000000;
		Dplus[4652] = 14'b0000000_0000000;
		Dplus[4653] = 14'b0000000_0000000;
		Dplus[4654] = 14'b0000000_0000000;
		Dplus[4655] = 14'b0000000_0000000;
		Dplus[4656] = 14'b0000000_0000000;
		Dplus[4657] = 14'b0000000_0000000;
		Dplus[4658] = 14'b0000000_0000000;
		Dplus[4659] = 14'b0000000_0000000;
		Dplus[4660] = 14'b0000000_0000000;
		Dplus[4661] = 14'b0000000_0000000;
		Dplus[4662] = 14'b0000000_0000000;
		Dplus[4663] = 14'b0000000_0000000;
		Dplus[4664] = 14'b0000000_0000000;
		Dplus[4665] = 14'b0000000_0000000;
		Dplus[4666] = 14'b0000000_0000000;
		Dplus[4667] = 14'b0000000_0000000;
		Dplus[4668] = 14'b0000000_0000000;
		Dplus[4669] = 14'b0000000_0000000;
		Dplus[4670] = 14'b0000000_0000000;
		Dplus[4671] = 14'b0000000_0000000;
		Dplus[4672] = 14'b0000000_0000000;
		Dplus[4673] = 14'b0000000_0000000;
		Dplus[4674] = 14'b0000000_0000000;
		Dplus[4675] = 14'b0000000_0000000;
		Dplus[4676] = 14'b0000000_0000000;
		Dplus[4677] = 14'b0000000_0000000;
		Dplus[4678] = 14'b0000000_0000000;
		Dplus[4679] = 14'b0000000_0000000;
		Dplus[4680] = 14'b0000000_0000000;
		Dplus[4681] = 14'b0000000_0000000;
		Dplus[4682] = 14'b0000000_0000000;
		Dplus[4683] = 14'b0000000_0000000;
		Dplus[4684] = 14'b0000000_0000000;
		Dplus[4685] = 14'b0000000_0000000;
		Dplus[4686] = 14'b0000000_0000000;
		Dplus[4687] = 14'b0000000_0000000;
		Dplus[4688] = 14'b0000000_0000000;
		Dplus[4689] = 14'b0000000_0000000;
		Dplus[4690] = 14'b0000000_0000000;
		Dplus[4691] = 14'b0000000_0000000;
		Dplus[4692] = 14'b0000000_0000000;
		Dplus[4693] = 14'b0000000_0000000;
		Dplus[4694] = 14'b0000000_0000000;
		Dplus[4695] = 14'b0000000_0000000;
		Dplus[4696] = 14'b0000000_0000000;
		Dplus[4697] = 14'b0000000_0000000;
		Dplus[4698] = 14'b0000000_0000000;
		Dplus[4699] = 14'b0000000_0000000;
		Dplus[4700] = 14'b0000000_0000000;
		Dplus[4701] = 14'b0000000_0000000;
		Dplus[4702] = 14'b0000000_0000000;
		Dplus[4703] = 14'b0000000_0000000;
		Dplus[4704] = 14'b0000000_0000000;
		Dplus[4705] = 14'b0000000_0000000;
		Dplus[4706] = 14'b0000000_0000000;
		Dplus[4707] = 14'b0000000_0000000;
		Dplus[4708] = 14'b0000000_0000000;
		Dplus[4709] = 14'b0000000_0000000;
		Dplus[4710] = 14'b0000000_0000000;
		Dplus[4711] = 14'b0000000_0000000;
		Dplus[4712] = 14'b0000000_0000000;
		Dplus[4713] = 14'b0000000_0000000;
		Dplus[4714] = 14'b0000000_0000000;
		Dplus[4715] = 14'b0000000_0000000;
		Dplus[4716] = 14'b0000000_0000000;
		Dplus[4717] = 14'b0000000_0000000;
		Dplus[4718] = 14'b0000000_0000000;
		Dplus[4719] = 14'b0000000_0000000;
		Dplus[4720] = 14'b0000000_0000000;
		Dplus[4721] = 14'b0000000_0000000;
		Dplus[4722] = 14'b0000000_0000000;
		Dplus[4723] = 14'b0000000_0000000;
		Dplus[4724] = 14'b0000000_0000000;
		Dplus[4725] = 14'b0000000_0000000;
		Dplus[4726] = 14'b0000000_0000000;
		Dplus[4727] = 14'b0000000_0000000;
		Dplus[4728] = 14'b0000000_0000000;
		Dplus[4729] = 14'b0000000_0000000;
		Dplus[4730] = 14'b0000000_0000000;
		Dplus[4731] = 14'b0000000_0000000;
		Dplus[4732] = 14'b0000000_0000000;
		Dplus[4733] = 14'b0000000_0000000;
		Dplus[4734] = 14'b0000000_0000000;
		Dplus[4735] = 14'b0000000_0000000;
		Dplus[4736] = 14'b0000000_0000000;
		Dplus[4737] = 14'b0000000_0000000;
		Dplus[4738] = 14'b0000000_0000000;
		Dplus[4739] = 14'b0000000_0000000;
		Dplus[4740] = 14'b0000000_0000000;
		Dplus[4741] = 14'b0000000_0000000;
		Dplus[4742] = 14'b0000000_0000000;
		Dplus[4743] = 14'b0000000_0000000;
		Dplus[4744] = 14'b0000000_0000000;
		Dplus[4745] = 14'b0000000_0000000;
		Dplus[4746] = 14'b0000000_0000000;
		Dplus[4747] = 14'b0000000_0000000;
		Dplus[4748] = 14'b0000000_0000000;
		Dplus[4749] = 14'b0000000_0000000;
		Dplus[4750] = 14'b0000000_0000000;
		Dplus[4751] = 14'b0000000_0000000;
		Dplus[4752] = 14'b0000000_0000000;
		Dplus[4753] = 14'b0000000_0000000;
		Dplus[4754] = 14'b0000000_0000000;
		Dplus[4755] = 14'b0000000_0000000;
		Dplus[4756] = 14'b0000000_0000000;
		Dplus[4757] = 14'b0000000_0000000;
		Dplus[4758] = 14'b0000000_0000000;
		Dplus[4759] = 14'b0000000_0000000;
		Dplus[4760] = 14'b0000000_0000000;
		Dplus[4761] = 14'b0000000_0000000;
		Dplus[4762] = 14'b0000000_0000000;
		Dplus[4763] = 14'b0000000_0000000;
		Dplus[4764] = 14'b0000000_0000000;
		Dplus[4765] = 14'b0000000_0000000;
		Dplus[4766] = 14'b0000000_0000000;
		Dplus[4767] = 14'b0000000_0000000;
		Dplus[4768] = 14'b0000000_0000000;
		Dplus[4769] = 14'b0000000_0000000;
		Dplus[4770] = 14'b0000000_0000000;
		Dplus[4771] = 14'b0000000_0000000;
		Dplus[4772] = 14'b0000000_0000000;
		Dplus[4773] = 14'b0000000_0000000;
		Dplus[4774] = 14'b0000000_0000000;
		Dplus[4775] = 14'b0000000_0000000;
		Dplus[4776] = 14'b0000000_0000000;
		Dplus[4777] = 14'b0000000_0000000;
		Dplus[4778] = 14'b0000000_0000000;
		Dplus[4779] = 14'b0000000_0000000;
		Dplus[4780] = 14'b0000000_0000000;
		Dplus[4781] = 14'b0000000_0000000;
		Dplus[4782] = 14'b0000000_0000000;
		Dplus[4783] = 14'b0000000_0000000;
		Dplus[4784] = 14'b0000000_0000000;
		Dplus[4785] = 14'b0000000_0000000;
		Dplus[4786] = 14'b0000000_0000000;
		Dplus[4787] = 14'b0000000_0000000;
		Dplus[4788] = 14'b0000000_0000000;
		Dplus[4789] = 14'b0000000_0000000;
		Dplus[4790] = 14'b0000000_0000000;
		Dplus[4791] = 14'b0000000_0000000;
		Dplus[4792] = 14'b0000000_0000000;
		Dplus[4793] = 14'b0000000_0000000;
		Dplus[4794] = 14'b0000000_0000000;
		Dplus[4795] = 14'b0000000_0000000;
		Dplus[4796] = 14'b0000000_0000000;
		Dplus[4797] = 14'b0000000_0000000;
		Dplus[4798] = 14'b0000000_0000000;
		Dplus[4799] = 14'b0000000_0000000;
		Dplus[4800] = 14'b0000000_0000000;
		Dplus[4801] = 14'b0000000_0000000;
		Dplus[4802] = 14'b0000000_0000000;
		Dplus[4803] = 14'b0000000_0000000;
		Dplus[4804] = 14'b0000000_0000000;
		Dplus[4805] = 14'b0000000_0000000;
		Dplus[4806] = 14'b0000000_0000000;
		Dplus[4807] = 14'b0000000_0000000;
		Dplus[4808] = 14'b0000000_0000000;
		Dplus[4809] = 14'b0000000_0000000;
		Dplus[4810] = 14'b0000000_0000000;
		Dplus[4811] = 14'b0000000_0000000;
		Dplus[4812] = 14'b0000000_0000000;
		Dplus[4813] = 14'b0000000_0000000;
		Dplus[4814] = 14'b0000000_0000000;
		Dplus[4815] = 14'b0000000_0000000;
		Dplus[4816] = 14'b0000000_0000000;
		Dplus[4817] = 14'b0000000_0000000;
		Dplus[4818] = 14'b0000000_0000000;
		Dplus[4819] = 14'b0000000_0000000;
		Dplus[4820] = 14'b0000000_0000000;
		Dplus[4821] = 14'b0000000_0000000;
		Dplus[4822] = 14'b0000000_0000000;
		Dplus[4823] = 14'b0000000_0000000;
		Dplus[4824] = 14'b0000000_0000000;
		Dplus[4825] = 14'b0000000_0000000;
		Dplus[4826] = 14'b0000000_0000000;
		Dplus[4827] = 14'b0000000_0000000;
		Dplus[4828] = 14'b0000000_0000000;
		Dplus[4829] = 14'b0000000_0000000;
		Dplus[4830] = 14'b0000000_0000000;
		Dplus[4831] = 14'b0000000_0000000;
		Dplus[4832] = 14'b0000000_0000000;
		Dplus[4833] = 14'b0000000_0000000;
		Dplus[4834] = 14'b0000000_0000000;
		Dplus[4835] = 14'b0000000_0000000;
		Dplus[4836] = 14'b0000000_0000000;
		Dplus[4837] = 14'b0000000_0000000;
		Dplus[4838] = 14'b0000000_0000000;
		Dplus[4839] = 14'b0000000_0000000;
		Dplus[4840] = 14'b0000000_0000000;
		Dplus[4841] = 14'b0000000_0000000;
		Dplus[4842] = 14'b0000000_0000000;
		Dplus[4843] = 14'b0000000_0000000;
		Dplus[4844] = 14'b0000000_0000000;
		Dplus[4845] = 14'b0000000_0000000;
		Dplus[4846] = 14'b0000000_0000000;
		Dplus[4847] = 14'b0000000_0000000;
		Dplus[4848] = 14'b0000000_0000000;
		Dplus[4849] = 14'b0000000_0000000;
		Dplus[4850] = 14'b0000000_0000000;
		Dplus[4851] = 14'b0000000_0000000;
		Dplus[4852] = 14'b0000000_0000000;
		Dplus[4853] = 14'b0000000_0000000;
		Dplus[4854] = 14'b0000000_0000000;
		Dplus[4855] = 14'b0000000_0000000;
		Dplus[4856] = 14'b0000000_0000000;
		Dplus[4857] = 14'b0000000_0000000;
		Dplus[4858] = 14'b0000000_0000000;
		Dplus[4859] = 14'b0000000_0000000;
		Dplus[4860] = 14'b0000000_0000000;
		Dplus[4861] = 14'b0000000_0000000;
		Dplus[4862] = 14'b0000000_0000000;
		Dplus[4863] = 14'b0000000_0000000;
		Dplus[4864] = 14'b0000000_0000000;
		Dplus[4865] = 14'b0000000_0000000;
		Dplus[4866] = 14'b0000000_0000000;
		Dplus[4867] = 14'b0000000_0000000;
		Dplus[4868] = 14'b0000000_0000000;
		Dplus[4869] = 14'b0000000_0000000;
		Dplus[4870] = 14'b0000000_0000000;
		Dplus[4871] = 14'b0000000_0000000;
		Dplus[4872] = 14'b0000000_0000000;
		Dplus[4873] = 14'b0000000_0000000;
		Dplus[4874] = 14'b0000000_0000000;
		Dplus[4875] = 14'b0000000_0000000;
		Dplus[4876] = 14'b0000000_0000000;
		Dplus[4877] = 14'b0000000_0000000;
		Dplus[4878] = 14'b0000000_0000000;
		Dplus[4879] = 14'b0000000_0000000;
		Dplus[4880] = 14'b0000000_0000000;
		Dplus[4881] = 14'b0000000_0000000;
		Dplus[4882] = 14'b0000000_0000000;
		Dplus[4883] = 14'b0000000_0000000;
		Dplus[4884] = 14'b0000000_0000000;
		Dplus[4885] = 14'b0000000_0000000;
		Dplus[4886] = 14'b0000000_0000000;
		Dplus[4887] = 14'b0000000_0000000;
		Dplus[4888] = 14'b0000000_0000000;
		Dplus[4889] = 14'b0000000_0000000;
		Dplus[4890] = 14'b0000000_0000000;
		Dplus[4891] = 14'b0000000_0000000;
		Dplus[4892] = 14'b0000000_0000000;
		Dplus[4893] = 14'b0000000_0000000;
		Dplus[4894] = 14'b0000000_0000000;
		Dplus[4895] = 14'b0000000_0000000;
		Dplus[4896] = 14'b0000000_0000000;
		Dplus[4897] = 14'b0000000_0000000;
		Dplus[4898] = 14'b0000000_0000000;
		Dplus[4899] = 14'b0000000_0000000;
		Dplus[4900] = 14'b0000000_0000000;
		Dplus[4901] = 14'b0000000_0000000;
		Dplus[4902] = 14'b0000000_0000000;
		Dplus[4903] = 14'b0000000_0000000;
		Dplus[4904] = 14'b0000000_0000000;
		Dplus[4905] = 14'b0000000_0000000;
		Dplus[4906] = 14'b0000000_0000000;
		Dplus[4907] = 14'b0000000_0000000;
		Dplus[4908] = 14'b0000000_0000000;
		Dplus[4909] = 14'b0000000_0000000;
		Dplus[4910] = 14'b0000000_0000000;
		Dplus[4911] = 14'b0000000_0000000;
		Dplus[4912] = 14'b0000000_0000000;
		Dplus[4913] = 14'b0000000_0000000;
		Dplus[4914] = 14'b0000000_0000000;
		Dplus[4915] = 14'b0000000_0000000;
		Dplus[4916] = 14'b0000000_0000000;
		Dplus[4917] = 14'b0000000_0000000;
		Dplus[4918] = 14'b0000000_0000000;
		Dplus[4919] = 14'b0000000_0000000;
		Dplus[4920] = 14'b0000000_0000000;
		Dplus[4921] = 14'b0000000_0000000;
		Dplus[4922] = 14'b0000000_0000000;
		Dplus[4923] = 14'b0000000_0000000;
		Dplus[4924] = 14'b0000000_0000000;
		Dplus[4925] = 14'b0000000_0000000;
		Dplus[4926] = 14'b0000000_0000000;
		Dplus[4927] = 14'b0000000_0000000;
		Dplus[4928] = 14'b0000000_0000000;
		Dplus[4929] = 14'b0000000_0000000;
		Dplus[4930] = 14'b0000000_0000000;
		Dplus[4931] = 14'b0000000_0000000;
		Dplus[4932] = 14'b0000000_0000000;
		Dplus[4933] = 14'b0000000_0000000;
		Dplus[4934] = 14'b0000000_0000000;
		Dplus[4935] = 14'b0000000_0000000;
		Dplus[4936] = 14'b0000000_0000000;
		Dplus[4937] = 14'b0000000_0000000;
		Dplus[4938] = 14'b0000000_0000000;
		Dplus[4939] = 14'b0000000_0000000;
		Dplus[4940] = 14'b0000000_0000000;
		Dplus[4941] = 14'b0000000_0000000;
		Dplus[4942] = 14'b0000000_0000000;
		Dplus[4943] = 14'b0000000_0000000;
		Dplus[4944] = 14'b0000000_0000000;
		Dplus[4945] = 14'b0000000_0000000;
		Dplus[4946] = 14'b0000000_0000000;
		Dplus[4947] = 14'b0000000_0000000;
		Dplus[4948] = 14'b0000000_0000000;
		Dplus[4949] = 14'b0000000_0000000;
		Dplus[4950] = 14'b0000000_0000000;
		Dplus[4951] = 14'b0000000_0000000;
		Dplus[4952] = 14'b0000000_0000000;
		Dplus[4953] = 14'b0000000_0000000;
		Dplus[4954] = 14'b0000000_0000000;
		Dplus[4955] = 14'b0000000_0000000;
		Dplus[4956] = 14'b0000000_0000000;
		Dplus[4957] = 14'b0000000_0000000;
		Dplus[4958] = 14'b0000000_0000000;
		Dplus[4959] = 14'b0000000_0000000;
		Dplus[4960] = 14'b0000000_0000000;
		Dplus[4961] = 14'b0000000_0000000;
		Dplus[4962] = 14'b0000000_0000000;
		Dplus[4963] = 14'b0000000_0000000;
		Dplus[4964] = 14'b0000000_0000000;
		Dplus[4965] = 14'b0000000_0000000;
		Dplus[4966] = 14'b0000000_0000000;
		Dplus[4967] = 14'b0000000_0000000;
		Dplus[4968] = 14'b0000000_0000000;
		Dplus[4969] = 14'b0000000_0000000;
		Dplus[4970] = 14'b0000000_0000000;
		Dplus[4971] = 14'b0000000_0000000;
		Dplus[4972] = 14'b0000000_0000000;
		Dplus[4973] = 14'b0000000_0000000;
		Dplus[4974] = 14'b0000000_0000000;
		Dplus[4975] = 14'b0000000_0000000;
		Dplus[4976] = 14'b0000000_0000000;
		Dplus[4977] = 14'b0000000_0000000;
		Dplus[4978] = 14'b0000000_0000000;
		Dplus[4979] = 14'b0000000_0000000;
		Dplus[4980] = 14'b0000000_0000000;
		Dplus[4981] = 14'b0000000_0000000;
		Dplus[4982] = 14'b0000000_0000000;
		Dplus[4983] = 14'b0000000_0000000;
		Dplus[4984] = 14'b0000000_0000000;
		Dplus[4985] = 14'b0000000_0000000;
		Dplus[4986] = 14'b0000000_0000000;
		Dplus[4987] = 14'b0000000_0000000;
		Dplus[4988] = 14'b0000000_0000000;
		Dplus[4989] = 14'b0000000_0000000;
		Dplus[4990] = 14'b0000000_0000000;
		Dplus[4991] = 14'b0000000_0000000;
		Dplus[4992] = 14'b0000000_0000000;
		Dplus[4993] = 14'b0000000_0000000;
		Dplus[4994] = 14'b0000000_0000000;
		Dplus[4995] = 14'b0000000_0000000;
		Dplus[4996] = 14'b0000000_0000000;
		Dplus[4997] = 14'b0000000_0000000;
		Dplus[4998] = 14'b0000000_0000000;
		Dplus[4999] = 14'b0000000_0000000;
		Dplus[5000] = 14'b0000000_0000000;
		Dplus[5001] = 14'b0000000_0000000;
		Dplus[5002] = 14'b0000000_0000000;
		Dplus[5003] = 14'b0000000_0000000;
		Dplus[5004] = 14'b0000000_0000000;
		Dplus[5005] = 14'b0000000_0000000;
		Dplus[5006] = 14'b0000000_0000000;
		Dplus[5007] = 14'b0000000_0000000;
		Dplus[5008] = 14'b0000000_0000000;
		Dplus[5009] = 14'b0000000_0000000;
		Dplus[5010] = 14'b0000000_0000000;
		Dplus[5011] = 14'b0000000_0000000;
		Dplus[5012] = 14'b0000000_0000000;
		Dplus[5013] = 14'b0000000_0000000;
		Dplus[5014] = 14'b0000000_0000000;
		Dplus[5015] = 14'b0000000_0000000;
		Dplus[5016] = 14'b0000000_0000000;
		Dplus[5017] = 14'b0000000_0000000;
		Dplus[5018] = 14'b0000000_0000000;
		Dplus[5019] = 14'b0000000_0000000;
		Dplus[5020] = 14'b0000000_0000000;
		Dplus[5021] = 14'b0000000_0000000;
		Dplus[5022] = 14'b0000000_0000000;
		Dplus[5023] = 14'b0000000_0000000;
		Dplus[5024] = 14'b0000000_0000000;
		Dplus[5025] = 14'b0000000_0000000;
		Dplus[5026] = 14'b0000000_0000000;
		Dplus[5027] = 14'b0000000_0000000;
		Dplus[5028] = 14'b0000000_0000000;
		Dplus[5029] = 14'b0000000_0000000;
		Dplus[5030] = 14'b0000000_0000000;
		Dplus[5031] = 14'b0000000_0000000;
		Dplus[5032] = 14'b0000000_0000000;
		Dplus[5033] = 14'b0000000_0000000;
		Dplus[5034] = 14'b0000000_0000000;
		Dplus[5035] = 14'b0000000_0000000;
		Dplus[5036] = 14'b0000000_0000000;
		Dplus[5037] = 14'b0000000_0000000;
		Dplus[5038] = 14'b0000000_0000000;
		Dplus[5039] = 14'b0000000_0000000;
		Dplus[5040] = 14'b0000000_0000000;
		Dplus[5041] = 14'b0000000_0000000;
		Dplus[5042] = 14'b0000000_0000000;
		Dplus[5043] = 14'b0000000_0000000;
		Dplus[5044] = 14'b0000000_0000000;
		Dplus[5045] = 14'b0000000_0000000;
		Dplus[5046] = 14'b0000000_0000000;
		Dplus[5047] = 14'b0000000_0000000;
		Dplus[5048] = 14'b0000000_0000000;
		Dplus[5049] = 14'b0000000_0000000;
		Dplus[5050] = 14'b0000000_0000000;
		Dplus[5051] = 14'b0000000_0000000;
		Dplus[5052] = 14'b0000000_0000000;
		Dplus[5053] = 14'b0000000_0000000;
		Dplus[5054] = 14'b0000000_0000000;
		Dplus[5055] = 14'b0000000_0000000;
		Dplus[5056] = 14'b0000000_0000000;
		Dplus[5057] = 14'b0000000_0000000;
		Dplus[5058] = 14'b0000000_0000000;
		Dplus[5059] = 14'b0000000_0000000;
		Dplus[5060] = 14'b0000000_0000000;
		Dplus[5061] = 14'b0000000_0000000;
		Dplus[5062] = 14'b0000000_0000000;
		Dplus[5063] = 14'b0000000_0000000;
		Dplus[5064] = 14'b0000000_0000000;
		Dplus[5065] = 14'b0000000_0000000;
		Dplus[5066] = 14'b0000000_0000000;
		Dplus[5067] = 14'b0000000_0000000;
		Dplus[5068] = 14'b0000000_0000000;
		Dplus[5069] = 14'b0000000_0000000;
		Dplus[5070] = 14'b0000000_0000000;
		Dplus[5071] = 14'b0000000_0000000;
		Dplus[5072] = 14'b0000000_0000000;
		Dplus[5073] = 14'b0000000_0000000;
		Dplus[5074] = 14'b0000000_0000000;
		Dplus[5075] = 14'b0000000_0000000;
		Dplus[5076] = 14'b0000000_0000000;
		Dplus[5077] = 14'b0000000_0000000;
		Dplus[5078] = 14'b0000000_0000000;
		Dplus[5079] = 14'b0000000_0000000;
		Dplus[5080] = 14'b0000000_0000000;
		Dplus[5081] = 14'b0000000_0000000;
		Dplus[5082] = 14'b0000000_0000000;
		Dplus[5083] = 14'b0000000_0000000;
		Dplus[5084] = 14'b0000000_0000000;
		Dplus[5085] = 14'b0000000_0000000;
		Dplus[5086] = 14'b0000000_0000000;
		Dplus[5087] = 14'b0000000_0000000;
		Dplus[5088] = 14'b0000000_0000000;
		Dplus[5089] = 14'b0000000_0000000;
		Dplus[5090] = 14'b0000000_0000000;
		Dplus[5091] = 14'b0000000_0000000;
		Dplus[5092] = 14'b0000000_0000000;
		Dplus[5093] = 14'b0000000_0000000;
		Dplus[5094] = 14'b0000000_0000000;
		Dplus[5095] = 14'b0000000_0000000;
		Dplus[5096] = 14'b0000000_0000000;
		Dplus[5097] = 14'b0000000_0000000;
		Dplus[5098] = 14'b0000000_0000000;
		Dplus[5099] = 14'b0000000_0000000;
		Dplus[5100] = 14'b0000000_0000000;
		Dplus[5101] = 14'b0000000_0000000;
		Dplus[5102] = 14'b0000000_0000000;
		Dplus[5103] = 14'b0000000_0000000;
		Dplus[5104] = 14'b0000000_0000000;
		Dplus[5105] = 14'b0000000_0000000;
		Dplus[5106] = 14'b0000000_0000000;
		Dplus[5107] = 14'b0000000_0000000;
		Dplus[5108] = 14'b0000000_0000000;
		Dplus[5109] = 14'b0000000_0000000;
		Dplus[5110] = 14'b0000000_0000000;
		Dplus[5111] = 14'b0000000_0000000;
		Dplus[5112] = 14'b0000000_0000000;
		Dplus[5113] = 14'b0000000_0000000;
		Dplus[5114] = 14'b0000000_0000000;
		Dplus[5115] = 14'b0000000_0000000;
		Dplus[5116] = 14'b0000000_0000000;
		Dplus[5117] = 14'b0000000_0000000;
		Dplus[5118] = 14'b0000000_0000000;
		Dplus[5119] = 14'b0000000_0000000;
		Dplus[5120] = 14'b0000000_0000000;
		Dplus[5121] = 14'b0000000_0000000;
		Dplus[5122] = 14'b0000000_0000000;
		Dplus[5123] = 14'b0000000_0000000;
		Dplus[5124] = 14'b0000000_0000000;
		Dplus[5125] = 14'b0000000_0000000;
		Dplus[5126] = 14'b0000000_0000000;
		Dplus[5127] = 14'b0000000_0000000;
		Dplus[5128] = 14'b0000000_0000000;
		Dplus[5129] = 14'b0000000_0000000;
		Dplus[5130] = 14'b0000000_0000000;
		Dplus[5131] = 14'b0000000_0000000;
		Dplus[5132] = 14'b0000000_0000000;
		Dplus[5133] = 14'b0000000_0000000;
		Dplus[5134] = 14'b0000000_0000000;
		Dplus[5135] = 14'b0000000_0000000;
		Dplus[5136] = 14'b0000000_0000000;
		Dplus[5137] = 14'b0000000_0000000;
		Dplus[5138] = 14'b0000000_0000000;
		Dplus[5139] = 14'b0000000_0000000;
		Dplus[5140] = 14'b0000000_0000000;
		Dplus[5141] = 14'b0000000_0000000;
		Dplus[5142] = 14'b0000000_0000000;
		Dplus[5143] = 14'b0000000_0000000;
		Dplus[5144] = 14'b0000000_0000000;
		Dplus[5145] = 14'b0000000_0000000;
		Dplus[5146] = 14'b0000000_0000000;
		Dplus[5147] = 14'b0000000_0000000;
		Dplus[5148] = 14'b0000000_0000000;
		Dplus[5149] = 14'b0000000_0000000;
		Dplus[5150] = 14'b0000000_0000000;
		Dplus[5151] = 14'b0000000_0000000;
		Dplus[5152] = 14'b0000000_0000000;
		Dplus[5153] = 14'b0000000_0000000;
		Dplus[5154] = 14'b0000000_0000000;
		Dplus[5155] = 14'b0000000_0000000;
		Dplus[5156] = 14'b0000000_0000000;
		Dplus[5157] = 14'b0000000_0000000;
		Dplus[5158] = 14'b0000000_0000000;
		Dplus[5159] = 14'b0000000_0000000;
		Dplus[5160] = 14'b0000000_0000000;
		Dplus[5161] = 14'b0000000_0000000;
		Dplus[5162] = 14'b0000000_0000000;
		Dplus[5163] = 14'b0000000_0000000;
		Dplus[5164] = 14'b0000000_0000000;
		Dplus[5165] = 14'b0000000_0000000;
		Dplus[5166] = 14'b0000000_0000000;
		Dplus[5167] = 14'b0000000_0000000;
		Dplus[5168] = 14'b0000000_0000000;
		Dplus[5169] = 14'b0000000_0000000;
		Dplus[5170] = 14'b0000000_0000000;
		Dplus[5171] = 14'b0000000_0000000;
		Dplus[5172] = 14'b0000000_0000000;
		Dplus[5173] = 14'b0000000_0000000;
		Dplus[5174] = 14'b0000000_0000000;
		Dplus[5175] = 14'b0000000_0000000;
		Dplus[5176] = 14'b0000000_0000000;
		Dplus[5177] = 14'b0000000_0000000;
		Dplus[5178] = 14'b0000000_0000000;
		Dplus[5179] = 14'b0000000_0000000;
		Dplus[5180] = 14'b0000000_0000000;
		Dplus[5181] = 14'b0000000_0000000;
		Dplus[5182] = 14'b0000000_0000000;
		Dplus[5183] = 14'b0000000_0000000;
		Dplus[5184] = 14'b0000000_0000000;
		Dplus[5185] = 14'b0000000_0000000;
		Dplus[5186] = 14'b0000000_0000000;
		Dplus[5187] = 14'b0000000_0000000;
		Dplus[5188] = 14'b0000000_0000000;
		Dplus[5189] = 14'b0000000_0000000;
		Dplus[5190] = 14'b0000000_0000000;
		Dplus[5191] = 14'b0000000_0000000;
		Dplus[5192] = 14'b0000000_0000000;
		Dplus[5193] = 14'b0000000_0000000;
		Dplus[5194] = 14'b0000000_0000000;
		Dplus[5195] = 14'b0000000_0000000;
		Dplus[5196] = 14'b0000000_0000000;
		Dplus[5197] = 14'b0000000_0000000;
		Dplus[5198] = 14'b0000000_0000000;
		Dplus[5199] = 14'b0000000_0000000;
		Dplus[5200] = 14'b0000000_0000000;
		Dplus[5201] = 14'b0000000_0000000;
		Dplus[5202] = 14'b0000000_0000000;
		Dplus[5203] = 14'b0000000_0000000;
		Dplus[5204] = 14'b0000000_0000000;
		Dplus[5205] = 14'b0000000_0000000;
		Dplus[5206] = 14'b0000000_0000000;
		Dplus[5207] = 14'b0000000_0000000;
		Dplus[5208] = 14'b0000000_0000000;
		Dplus[5209] = 14'b0000000_0000000;
		Dplus[5210] = 14'b0000000_0000000;
		Dplus[5211] = 14'b0000000_0000000;
		Dplus[5212] = 14'b0000000_0000000;
		Dplus[5213] = 14'b0000000_0000000;
		Dplus[5214] = 14'b0000000_0000000;
		Dplus[5215] = 14'b0000000_0000000;
		Dplus[5216] = 14'b0000000_0000000;
		Dplus[5217] = 14'b0000000_0000000;
		Dplus[5218] = 14'b0000000_0000000;
		Dplus[5219] = 14'b0000000_0000000;
		Dplus[5220] = 14'b0000000_0000000;
		Dplus[5221] = 14'b0000000_0000000;
		Dplus[5222] = 14'b0000000_0000000;
		Dplus[5223] = 14'b0000000_0000000;
		Dplus[5224] = 14'b0000000_0000000;
		Dplus[5225] = 14'b0000000_0000000;
		Dplus[5226] = 14'b0000000_0000000;
		Dplus[5227] = 14'b0000000_0000000;
		Dplus[5228] = 14'b0000000_0000000;
		Dplus[5229] = 14'b0000000_0000000;
		Dplus[5230] = 14'b0000000_0000000;
		Dplus[5231] = 14'b0000000_0000000;
		Dplus[5232] = 14'b0000000_0000000;
		Dplus[5233] = 14'b0000000_0000000;
		Dplus[5234] = 14'b0000000_0000000;
		Dplus[5235] = 14'b0000000_0000000;
		Dplus[5236] = 14'b0000000_0000000;
		Dplus[5237] = 14'b0000000_0000000;
		Dplus[5238] = 14'b0000000_0000000;
		Dplus[5239] = 14'b0000000_0000000;
		Dplus[5240] = 14'b0000000_0000000;
		Dplus[5241] = 14'b0000000_0000000;
		Dplus[5242] = 14'b0000000_0000000;
		Dplus[5243] = 14'b0000000_0000000;
		Dplus[5244] = 14'b0000000_0000000;
		Dplus[5245] = 14'b0000000_0000000;
		Dplus[5246] = 14'b0000000_0000000;
		Dplus[5247] = 14'b0000000_0000000;
		Dplus[5248] = 14'b0000000_0000000;
		Dplus[5249] = 14'b0000000_0000000;
		Dplus[5250] = 14'b0000000_0000000;
		Dplus[5251] = 14'b0000000_0000000;
		Dplus[5252] = 14'b0000000_0000000;
		Dplus[5253] = 14'b0000000_0000000;
		Dplus[5254] = 14'b0000000_0000000;
		Dplus[5255] = 14'b0000000_0000000;
		Dplus[5256] = 14'b0000000_0000000;
		Dplus[5257] = 14'b0000000_0000000;
		Dplus[5258] = 14'b0000000_0000000;
		Dplus[5259] = 14'b0000000_0000000;
		Dplus[5260] = 14'b0000000_0000000;
		Dplus[5261] = 14'b0000000_0000000;
		Dplus[5262] = 14'b0000000_0000000;
		Dplus[5263] = 14'b0000000_0000000;
		Dplus[5264] = 14'b0000000_0000000;
		Dplus[5265] = 14'b0000000_0000000;
		Dplus[5266] = 14'b0000000_0000000;
		Dplus[5267] = 14'b0000000_0000000;
		Dplus[5268] = 14'b0000000_0000000;
		Dplus[5269] = 14'b0000000_0000000;
		Dplus[5270] = 14'b0000000_0000000;
		Dplus[5271] = 14'b0000000_0000000;
		Dplus[5272] = 14'b0000000_0000000;
		Dplus[5273] = 14'b0000000_0000000;
		Dplus[5274] = 14'b0000000_0000000;
		Dplus[5275] = 14'b0000000_0000000;
		Dplus[5276] = 14'b0000000_0000000;
		Dplus[5277] = 14'b0000000_0000000;
		Dplus[5278] = 14'b0000000_0000000;
		Dplus[5279] = 14'b0000000_0000000;
		Dplus[5280] = 14'b0000000_0000000;
		Dplus[5281] = 14'b0000000_0000000;
		Dplus[5282] = 14'b0000000_0000000;
		Dplus[5283] = 14'b0000000_0000000;
		Dplus[5284] = 14'b0000000_0000000;
		Dplus[5285] = 14'b0000000_0000000;
		Dplus[5286] = 14'b0000000_0000000;
		Dplus[5287] = 14'b0000000_0000000;
		Dplus[5288] = 14'b0000000_0000000;
		Dplus[5289] = 14'b0000000_0000000;
		Dplus[5290] = 14'b0000000_0000000;
		Dplus[5291] = 14'b0000000_0000000;
		Dplus[5292] = 14'b0000000_0000000;
		Dplus[5293] = 14'b0000000_0000000;
		Dplus[5294] = 14'b0000000_0000000;
		Dplus[5295] = 14'b0000000_0000000;
		Dplus[5296] = 14'b0000000_0000000;
		Dplus[5297] = 14'b0000000_0000000;
		Dplus[5298] = 14'b0000000_0000000;
		Dplus[5299] = 14'b0000000_0000000;
		Dplus[5300] = 14'b0000000_0000000;
		Dplus[5301] = 14'b0000000_0000000;
		Dplus[5302] = 14'b0000000_0000000;
		Dplus[5303] = 14'b0000000_0000000;
		Dplus[5304] = 14'b0000000_0000000;
		Dplus[5305] = 14'b0000000_0000000;
		Dplus[5306] = 14'b0000000_0000000;
		Dplus[5307] = 14'b0000000_0000000;
		Dplus[5308] = 14'b0000000_0000000;
		Dplus[5309] = 14'b0000000_0000000;
		Dplus[5310] = 14'b0000000_0000000;
		Dplus[5311] = 14'b0000000_0000000;
		Dplus[5312] = 14'b0000000_0000000;
		Dplus[5313] = 14'b0000000_0000000;
		Dplus[5314] = 14'b0000000_0000000;
		Dplus[5315] = 14'b0000000_0000000;
		Dplus[5316] = 14'b0000000_0000000;
		Dplus[5317] = 14'b0000000_0000000;
		Dplus[5318] = 14'b0000000_0000000;
		Dplus[5319] = 14'b0000000_0000000;
		Dplus[5320] = 14'b0000000_0000000;
		Dplus[5321] = 14'b0000000_0000000;
		Dplus[5322] = 14'b0000000_0000000;
		Dplus[5323] = 14'b0000000_0000000;
		Dplus[5324] = 14'b0000000_0000000;
		Dplus[5325] = 14'b0000000_0000000;
		Dplus[5326] = 14'b0000000_0000000;
		Dplus[5327] = 14'b0000000_0000000;
		Dplus[5328] = 14'b0000000_0000000;
		Dplus[5329] = 14'b0000000_0000000;
		Dplus[5330] = 14'b0000000_0000000;
		Dplus[5331] = 14'b0000000_0000000;
		Dplus[5332] = 14'b0000000_0000000;
		Dplus[5333] = 14'b0000000_0000000;
		Dplus[5334] = 14'b0000000_0000000;
		Dplus[5335] = 14'b0000000_0000000;
		Dplus[5336] = 14'b0000000_0000000;
		Dplus[5337] = 14'b0000000_0000000;
		Dplus[5338] = 14'b0000000_0000000;
		Dplus[5339] = 14'b0000000_0000000;
		Dplus[5340] = 14'b0000000_0000000;
		Dplus[5341] = 14'b0000000_0000000;
		Dplus[5342] = 14'b0000000_0000000;
		Dplus[5343] = 14'b0000000_0000000;
		Dplus[5344] = 14'b0000000_0000000;
		Dplus[5345] = 14'b0000000_0000000;
		Dplus[5346] = 14'b0000000_0000000;
		Dplus[5347] = 14'b0000000_0000000;
		Dplus[5348] = 14'b0000000_0000000;
		Dplus[5349] = 14'b0000000_0000000;
		Dplus[5350] = 14'b0000000_0000000;
		Dplus[5351] = 14'b0000000_0000000;
		Dplus[5352] = 14'b0000000_0000000;
		Dplus[5353] = 14'b0000000_0000000;
		Dplus[5354] = 14'b0000000_0000000;
		Dplus[5355] = 14'b0000000_0000000;
		Dplus[5356] = 14'b0000000_0000000;
		Dplus[5357] = 14'b0000000_0000000;
		Dplus[5358] = 14'b0000000_0000000;
		Dplus[5359] = 14'b0000000_0000000;
		Dplus[5360] = 14'b0000000_0000000;
		Dplus[5361] = 14'b0000000_0000000;
		Dplus[5362] = 14'b0000000_0000000;
		Dplus[5363] = 14'b0000000_0000000;
		Dplus[5364] = 14'b0000000_0000000;
		Dplus[5365] = 14'b0000000_0000000;
		Dplus[5366] = 14'b0000000_0000000;
		Dplus[5367] = 14'b0000000_0000000;
		Dplus[5368] = 14'b0000000_0000000;
		Dplus[5369] = 14'b0000000_0000000;
		Dplus[5370] = 14'b0000000_0000000;
		Dplus[5371] = 14'b0000000_0000000;
		Dplus[5372] = 14'b0000000_0000000;
		Dplus[5373] = 14'b0000000_0000000;
		Dplus[5374] = 14'b0000000_0000000;
		Dplus[5375] = 14'b0000000_0000000;
		Dplus[5376] = 14'b0000000_0000000;
		Dplus[5377] = 14'b0000000_0000000;
		Dplus[5378] = 14'b0000000_0000000;
		Dplus[5379] = 14'b0000000_0000000;
		Dplus[5380] = 14'b0000000_0000000;
		Dplus[5381] = 14'b0000000_0000000;
		Dplus[5382] = 14'b0000000_0000000;
		Dplus[5383] = 14'b0000000_0000000;
		Dplus[5384] = 14'b0000000_0000000;
		Dplus[5385] = 14'b0000000_0000000;
		Dplus[5386] = 14'b0000000_0000000;
		Dplus[5387] = 14'b0000000_0000000;
		Dplus[5388] = 14'b0000000_0000000;
		Dplus[5389] = 14'b0000000_0000000;
		Dplus[5390] = 14'b0000000_0000000;
		Dplus[5391] = 14'b0000000_0000000;
		Dplus[5392] = 14'b0000000_0000000;
		Dplus[5393] = 14'b0000000_0000000;
		Dplus[5394] = 14'b0000000_0000000;
		Dplus[5395] = 14'b0000000_0000000;
		Dplus[5396] = 14'b0000000_0000000;
		Dplus[5397] = 14'b0000000_0000000;
		Dplus[5398] = 14'b0000000_0000000;
		Dplus[5399] = 14'b0000000_0000000;
		Dplus[5400] = 14'b0000000_0000000;
		Dplus[5401] = 14'b0000000_0000000;
		Dplus[5402] = 14'b0000000_0000000;
		Dplus[5403] = 14'b0000000_0000000;
		Dplus[5404] = 14'b0000000_0000000;
		Dplus[5405] = 14'b0000000_0000000;
		Dplus[5406] = 14'b0000000_0000000;
		Dplus[5407] = 14'b0000000_0000000;
		Dplus[5408] = 14'b0000000_0000000;
		Dplus[5409] = 14'b0000000_0000000;
		Dplus[5410] = 14'b0000000_0000000;
		Dplus[5411] = 14'b0000000_0000000;
		Dplus[5412] = 14'b0000000_0000000;
		Dplus[5413] = 14'b0000000_0000000;
		Dplus[5414] = 14'b0000000_0000000;
		Dplus[5415] = 14'b0000000_0000000;
		Dplus[5416] = 14'b0000000_0000000;
		Dplus[5417] = 14'b0000000_0000000;
		Dplus[5418] = 14'b0000000_0000000;
		Dplus[5419] = 14'b0000000_0000000;
		Dplus[5420] = 14'b0000000_0000000;
		Dplus[5421] = 14'b0000000_0000000;
		Dplus[5422] = 14'b0000000_0000000;
		Dplus[5423] = 14'b0000000_0000000;
		Dplus[5424] = 14'b0000000_0000000;
		Dplus[5425] = 14'b0000000_0000000;
		Dplus[5426] = 14'b0000000_0000000;
		Dplus[5427] = 14'b0000000_0000000;
		Dplus[5428] = 14'b0000000_0000000;
		Dplus[5429] = 14'b0000000_0000000;
		Dplus[5430] = 14'b0000000_0000000;
		Dplus[5431] = 14'b0000000_0000000;
		Dplus[5432] = 14'b0000000_0000000;
		Dplus[5433] = 14'b0000000_0000000;
		Dplus[5434] = 14'b0000000_0000000;
		Dplus[5435] = 14'b0000000_0000000;
		Dplus[5436] = 14'b0000000_0000000;
		Dplus[5437] = 14'b0000000_0000000;
		Dplus[5438] = 14'b0000000_0000000;
		Dplus[5439] = 14'b0000000_0000000;
		Dplus[5440] = 14'b0000000_0000000;
		Dplus[5441] = 14'b0000000_0000000;
		Dplus[5442] = 14'b0000000_0000000;
		Dplus[5443] = 14'b0000000_0000000;
		Dplus[5444] = 14'b0000000_0000000;
		Dplus[5445] = 14'b0000000_0000000;
		Dplus[5446] = 14'b0000000_0000000;
		Dplus[5447] = 14'b0000000_0000000;
		Dplus[5448] = 14'b0000000_0000000;
		Dplus[5449] = 14'b0000000_0000000;
		Dplus[5450] = 14'b0000000_0000000;
		Dplus[5451] = 14'b0000000_0000000;
		Dplus[5452] = 14'b0000000_0000000;
		Dplus[5453] = 14'b0000000_0000000;
		Dplus[5454] = 14'b0000000_0000000;
		Dplus[5455] = 14'b0000000_0000000;
		Dplus[5456] = 14'b0000000_0000000;
		Dplus[5457] = 14'b0000000_0000000;
		Dplus[5458] = 14'b0000000_0000000;
		Dplus[5459] = 14'b0000000_0000000;
		Dplus[5460] = 14'b0000000_0000000;
		Dplus[5461] = 14'b0000000_0000000;
		Dplus[5462] = 14'b0000000_0000000;
		Dplus[5463] = 14'b0000000_0000000;
		Dplus[5464] = 14'b0000000_0000000;
		Dplus[5465] = 14'b0000000_0000000;
		Dplus[5466] = 14'b0000000_0000000;
		Dplus[5467] = 14'b0000000_0000000;
		Dplus[5468] = 14'b0000000_0000000;
		Dplus[5469] = 14'b0000000_0000000;
		Dplus[5470] = 14'b0000000_0000000;
		Dplus[5471] = 14'b0000000_0000000;
		Dplus[5472] = 14'b0000000_0000000;
		Dplus[5473] = 14'b0000000_0000000;
		Dplus[5474] = 14'b0000000_0000000;
		Dplus[5475] = 14'b0000000_0000000;
		Dplus[5476] = 14'b0000000_0000000;
		Dplus[5477] = 14'b0000000_0000000;
		Dplus[5478] = 14'b0000000_0000000;
		Dplus[5479] = 14'b0000000_0000000;
		Dplus[5480] = 14'b0000000_0000000;
		Dplus[5481] = 14'b0000000_0000000;
		Dplus[5482] = 14'b0000000_0000000;
		Dplus[5483] = 14'b0000000_0000000;
		Dplus[5484] = 14'b0000000_0000000;
		Dplus[5485] = 14'b0000000_0000000;
		Dplus[5486] = 14'b0000000_0000000;
		Dplus[5487] = 14'b0000000_0000000;
		Dplus[5488] = 14'b0000000_0000000;
		Dplus[5489] = 14'b0000000_0000000;
		Dplus[5490] = 14'b0000000_0000000;
		Dplus[5491] = 14'b0000000_0000000;
		Dplus[5492] = 14'b0000000_0000000;
		Dplus[5493] = 14'b0000000_0000000;
		Dplus[5494] = 14'b0000000_0000000;
		Dplus[5495] = 14'b0000000_0000000;
		Dplus[5496] = 14'b0000000_0000000;
		Dplus[5497] = 14'b0000000_0000000;
		Dplus[5498] = 14'b0000000_0000000;
		Dplus[5499] = 14'b0000000_0000000;
		Dplus[5500] = 14'b0000000_0000000;
		Dplus[5501] = 14'b0000000_0000000;
		Dplus[5502] = 14'b0000000_0000000;
		Dplus[5503] = 14'b0000000_0000000;
		Dplus[5504] = 14'b0000000_0000000;
		Dplus[5505] = 14'b0000000_0000000;
		Dplus[5506] = 14'b0000000_0000000;
		Dplus[5507] = 14'b0000000_0000000;
		Dplus[5508] = 14'b0000000_0000000;
		Dplus[5509] = 14'b0000000_0000000;
		Dplus[5510] = 14'b0000000_0000000;
		Dplus[5511] = 14'b0000000_0000000;
		Dplus[5512] = 14'b0000000_0000000;
		Dplus[5513] = 14'b0000000_0000000;
		Dplus[5514] = 14'b0000000_0000000;
		Dplus[5515] = 14'b0000000_0000000;
		Dplus[5516] = 14'b0000000_0000000;
		Dplus[5517] = 14'b0000000_0000000;
		Dplus[5518] = 14'b0000000_0000000;
		Dplus[5519] = 14'b0000000_0000000;
		Dplus[5520] = 14'b0000000_0000000;
		Dplus[5521] = 14'b0000000_0000000;
		Dplus[5522] = 14'b0000000_0000000;
		Dplus[5523] = 14'b0000000_0000000;
		Dplus[5524] = 14'b0000000_0000000;
		Dplus[5525] = 14'b0000000_0000000;
		Dplus[5526] = 14'b0000000_0000000;
		Dplus[5527] = 14'b0000000_0000000;
		Dplus[5528] = 14'b0000000_0000000;
		Dplus[5529] = 14'b0000000_0000000;
		Dplus[5530] = 14'b0000000_0000000;
		Dplus[5531] = 14'b0000000_0000000;
		Dplus[5532] = 14'b0000000_0000000;
		Dplus[5533] = 14'b0000000_0000000;
		Dplus[5534] = 14'b0000000_0000000;
		Dplus[5535] = 14'b0000000_0000000;
		Dplus[5536] = 14'b0000000_0000000;
		Dplus[5537] = 14'b0000000_0000000;
		Dplus[5538] = 14'b0000000_0000000;
		Dplus[5539] = 14'b0000000_0000000;
		Dplus[5540] = 14'b0000000_0000000;
		Dplus[5541] = 14'b0000000_0000000;
		Dplus[5542] = 14'b0000000_0000000;
		Dplus[5543] = 14'b0000000_0000000;
		Dplus[5544] = 14'b0000000_0000000;
		Dplus[5545] = 14'b0000000_0000000;
		Dplus[5546] = 14'b0000000_0000000;
		Dplus[5547] = 14'b0000000_0000000;
		Dplus[5548] = 14'b0000000_0000000;
		Dplus[5549] = 14'b0000000_0000000;
		Dplus[5550] = 14'b0000000_0000000;
		Dplus[5551] = 14'b0000000_0000000;
		Dplus[5552] = 14'b0000000_0000000;
		Dplus[5553] = 14'b0000000_0000000;
		Dplus[5554] = 14'b0000000_0000000;
		Dplus[5555] = 14'b0000000_0000000;
		Dplus[5556] = 14'b0000000_0000000;
		Dplus[5557] = 14'b0000000_0000000;
		Dplus[5558] = 14'b0000000_0000000;
		Dplus[5559] = 14'b0000000_0000000;
		Dplus[5560] = 14'b0000000_0000000;
		Dplus[5561] = 14'b0000000_0000000;
		Dplus[5562] = 14'b0000000_0000000;
		Dplus[5563] = 14'b0000000_0000000;
		Dplus[5564] = 14'b0000000_0000000;
		Dplus[5565] = 14'b0000000_0000000;
		Dplus[5566] = 14'b0000000_0000000;
		Dplus[5567] = 14'b0000000_0000000;
		Dplus[5568] = 14'b0000000_0000000;
		Dplus[5569] = 14'b0000000_0000000;
		Dplus[5570] = 14'b0000000_0000000;
		Dplus[5571] = 14'b0000000_0000000;
		Dplus[5572] = 14'b0000000_0000000;
		Dplus[5573] = 14'b0000000_0000000;
		Dplus[5574] = 14'b0000000_0000000;
		Dplus[5575] = 14'b0000000_0000000;
		Dplus[5576] = 14'b0000000_0000000;
		Dplus[5577] = 14'b0000000_0000000;
		Dplus[5578] = 14'b0000000_0000000;
		Dplus[5579] = 14'b0000000_0000000;
		Dplus[5580] = 14'b0000000_0000000;
		Dplus[5581] = 14'b0000000_0000000;
		Dplus[5582] = 14'b0000000_0000000;
		Dplus[5583] = 14'b0000000_0000000;
		Dplus[5584] = 14'b0000000_0000000;
		Dplus[5585] = 14'b0000000_0000000;
		Dplus[5586] = 14'b0000000_0000000;
		Dplus[5587] = 14'b0000000_0000000;
		Dplus[5588] = 14'b0000000_0000000;
		Dplus[5589] = 14'b0000000_0000000;
		Dplus[5590] = 14'b0000000_0000000;
		Dplus[5591] = 14'b0000000_0000000;
		Dplus[5592] = 14'b0000000_0000000;
		Dplus[5593] = 14'b0000000_0000000;
		Dplus[5594] = 14'b0000000_0000000;
		Dplus[5595] = 14'b0000000_0000000;
		Dplus[5596] = 14'b0000000_0000000;
		Dplus[5597] = 14'b0000000_0000000;
		Dplus[5598] = 14'b0000000_0000000;
		Dplus[5599] = 14'b0000000_0000000;
		Dplus[5600] = 14'b0000000_0000000;
		Dplus[5601] = 14'b0000000_0000000;
		Dplus[5602] = 14'b0000000_0000000;
		Dplus[5603] = 14'b0000000_0000000;
		Dplus[5604] = 14'b0000000_0000000;
		Dplus[5605] = 14'b0000000_0000000;
		Dplus[5606] = 14'b0000000_0000000;
		Dplus[5607] = 14'b0000000_0000000;
		Dplus[5608] = 14'b0000000_0000000;
		Dplus[5609] = 14'b0000000_0000000;
		Dplus[5610] = 14'b0000000_0000000;
		Dplus[5611] = 14'b0000000_0000000;
		Dplus[5612] = 14'b0000000_0000000;
		Dplus[5613] = 14'b0000000_0000000;
		Dplus[5614] = 14'b0000000_0000000;
		Dplus[5615] = 14'b0000000_0000000;
		Dplus[5616] = 14'b0000000_0000000;
		Dplus[5617] = 14'b0000000_0000000;
		Dplus[5618] = 14'b0000000_0000000;
		Dplus[5619] = 14'b0000000_0000000;
		Dplus[5620] = 14'b0000000_0000000;
		Dplus[5621] = 14'b0000000_0000000;
		Dplus[5622] = 14'b0000000_0000000;
		Dplus[5623] = 14'b0000000_0000000;
		Dplus[5624] = 14'b0000000_0000000;
		Dplus[5625] = 14'b0000000_0000000;
		Dplus[5626] = 14'b0000000_0000000;
		Dplus[5627] = 14'b0000000_0000000;
		Dplus[5628] = 14'b0000000_0000000;
		Dplus[5629] = 14'b0000000_0000000;
		Dplus[5630] = 14'b0000000_0000000;
		Dplus[5631] = 14'b0000000_0000000;
		Dplus[5632] = 14'b0000000_0000000;
		Dplus[5633] = 14'b0000000_0000000;
		Dplus[5634] = 14'b0000000_0000000;
		Dplus[5635] = 14'b0000000_0000000;
		Dplus[5636] = 14'b0000000_0000000;
		Dplus[5637] = 14'b0000000_0000000;
		Dplus[5638] = 14'b0000000_0000000;
		Dplus[5639] = 14'b0000000_0000000;
		Dplus[5640] = 14'b0000000_0000000;
		Dplus[5641] = 14'b0000000_0000000;
		Dplus[5642] = 14'b0000000_0000000;
		Dplus[5643] = 14'b0000000_0000000;
		Dplus[5644] = 14'b0000000_0000000;
		Dplus[5645] = 14'b0000000_0000000;
		Dplus[5646] = 14'b0000000_0000000;
		Dplus[5647] = 14'b0000000_0000000;
		Dplus[5648] = 14'b0000000_0000000;
		Dplus[5649] = 14'b0000000_0000000;
		Dplus[5650] = 14'b0000000_0000000;
		Dplus[5651] = 14'b0000000_0000000;
		Dplus[5652] = 14'b0000000_0000000;
		Dplus[5653] = 14'b0000000_0000000;
		Dplus[5654] = 14'b0000000_0000000;
		Dplus[5655] = 14'b0000000_0000000;
		Dplus[5656] = 14'b0000000_0000000;
		Dplus[5657] = 14'b0000000_0000000;
		Dplus[5658] = 14'b0000000_0000000;
		Dplus[5659] = 14'b0000000_0000000;
		Dplus[5660] = 14'b0000000_0000000;
		Dplus[5661] = 14'b0000000_0000000;
		Dplus[5662] = 14'b0000000_0000000;
		Dplus[5663] = 14'b0000000_0000000;
		Dplus[5664] = 14'b0000000_0000000;
		Dplus[5665] = 14'b0000000_0000000;
		Dplus[5666] = 14'b0000000_0000000;
		Dplus[5667] = 14'b0000000_0000000;
		Dplus[5668] = 14'b0000000_0000000;
		Dplus[5669] = 14'b0000000_0000000;
		Dplus[5670] = 14'b0000000_0000000;
		Dplus[5671] = 14'b0000000_0000000;
		Dplus[5672] = 14'b0000000_0000000;
		Dplus[5673] = 14'b0000000_0000000;
		Dplus[5674] = 14'b0000000_0000000;
		Dplus[5675] = 14'b0000000_0000000;
		Dplus[5676] = 14'b0000000_0000000;
		Dplus[5677] = 14'b0000000_0000000;
		Dplus[5678] = 14'b0000000_0000000;
		Dplus[5679] = 14'b0000000_0000000;
		Dplus[5680] = 14'b0000000_0000000;
		Dplus[5681] = 14'b0000000_0000000;
		Dplus[5682] = 14'b0000000_0000000;
		Dplus[5683] = 14'b0000000_0000000;
		Dplus[5684] = 14'b0000000_0000000;
		Dplus[5685] = 14'b0000000_0000000;
		Dplus[5686] = 14'b0000000_0000000;
		Dplus[5687] = 14'b0000000_0000000;
		Dplus[5688] = 14'b0000000_0000000;
		Dplus[5689] = 14'b0000000_0000000;
		Dplus[5690] = 14'b0000000_0000000;
		Dplus[5691] = 14'b0000000_0000000;
		Dplus[5692] = 14'b0000000_0000000;
		Dplus[5693] = 14'b0000000_0000000;
		Dplus[5694] = 14'b0000000_0000000;
		Dplus[5695] = 14'b0000000_0000000;
		Dplus[5696] = 14'b0000000_0000000;
		Dplus[5697] = 14'b0000000_0000000;
		Dplus[5698] = 14'b0000000_0000000;
		Dplus[5699] = 14'b0000000_0000000;
		Dplus[5700] = 14'b0000000_0000000;
		Dplus[5701] = 14'b0000000_0000000;
		Dplus[5702] = 14'b0000000_0000000;
		Dplus[5703] = 14'b0000000_0000000;
		Dplus[5704] = 14'b0000000_0000000;
		Dplus[5705] = 14'b0000000_0000000;
		Dplus[5706] = 14'b0000000_0000000;
		Dplus[5707] = 14'b0000000_0000000;
		Dplus[5708] = 14'b0000000_0000000;
		Dplus[5709] = 14'b0000000_0000000;
		Dplus[5710] = 14'b0000000_0000000;
		Dplus[5711] = 14'b0000000_0000000;
		Dplus[5712] = 14'b0000000_0000000;
		Dplus[5713] = 14'b0000000_0000000;
		Dplus[5714] = 14'b0000000_0000000;
		Dplus[5715] = 14'b0000000_0000000;
		Dplus[5716] = 14'b0000000_0000000;
		Dplus[5717] = 14'b0000000_0000000;
		Dplus[5718] = 14'b0000000_0000000;
		Dplus[5719] = 14'b0000000_0000000;
		Dplus[5720] = 14'b0000000_0000000;
		Dplus[5721] = 14'b0000000_0000000;
		Dplus[5722] = 14'b0000000_0000000;
		Dplus[5723] = 14'b0000000_0000000;
		Dplus[5724] = 14'b0000000_0000000;
		Dplus[5725] = 14'b0000000_0000000;
		Dplus[5726] = 14'b0000000_0000000;
		Dplus[5727] = 14'b0000000_0000000;
		Dplus[5728] = 14'b0000000_0000000;
		Dplus[5729] = 14'b0000000_0000000;
		Dplus[5730] = 14'b0000000_0000000;
		Dplus[5731] = 14'b0000000_0000000;
		Dplus[5732] = 14'b0000000_0000000;
		Dplus[5733] = 14'b0000000_0000000;
		Dplus[5734] = 14'b0000000_0000000;
		Dplus[5735] = 14'b0000000_0000000;
		Dplus[5736] = 14'b0000000_0000000;
		Dplus[5737] = 14'b0000000_0000000;
		Dplus[5738] = 14'b0000000_0000000;
		Dplus[5739] = 14'b0000000_0000000;
		Dplus[5740] = 14'b0000000_0000000;
		Dplus[5741] = 14'b0000000_0000000;
		Dplus[5742] = 14'b0000000_0000000;
		Dplus[5743] = 14'b0000000_0000000;
		Dplus[5744] = 14'b0000000_0000000;
		Dplus[5745] = 14'b0000000_0000000;
		Dplus[5746] = 14'b0000000_0000000;
		Dplus[5747] = 14'b0000000_0000000;
		Dplus[5748] = 14'b0000000_0000000;
		Dplus[5749] = 14'b0000000_0000000;
		Dplus[5750] = 14'b0000000_0000000;
		Dplus[5751] = 14'b0000000_0000000;
		Dplus[5752] = 14'b0000000_0000000;
		Dplus[5753] = 14'b0000000_0000000;
		Dplus[5754] = 14'b0000000_0000000;
		Dplus[5755] = 14'b0000000_0000000;
		Dplus[5756] = 14'b0000000_0000000;
		Dplus[5757] = 14'b0000000_0000000;
		Dplus[5758] = 14'b0000000_0000000;
		Dplus[5759] = 14'b0000000_0000000;
		Dplus[5760] = 14'b0000000_0000000;
		Dplus[5761] = 14'b0000000_0000000;
		Dplus[5762] = 14'b0000000_0000000;
		Dplus[5763] = 14'b0000000_0000000;
		Dplus[5764] = 14'b0000000_0000000;
		Dplus[5765] = 14'b0000000_0000000;
		Dplus[5766] = 14'b0000000_0000000;
		Dplus[5767] = 14'b0000000_0000000;
		Dplus[5768] = 14'b0000000_0000000;
		Dplus[5769] = 14'b0000000_0000000;
		Dplus[5770] = 14'b0000000_0000000;
		Dplus[5771] = 14'b0000000_0000000;
		Dplus[5772] = 14'b0000000_0000000;
		Dplus[5773] = 14'b0000000_0000000;
		Dplus[5774] = 14'b0000000_0000000;
		Dplus[5775] = 14'b0000000_0000000;
		Dplus[5776] = 14'b0000000_0000000;
		Dplus[5777] = 14'b0000000_0000000;
		Dplus[5778] = 14'b0000000_0000000;
		Dplus[5779] = 14'b0000000_0000000;
		Dplus[5780] = 14'b0000000_0000000;
		Dplus[5781] = 14'b0000000_0000000;
		Dplus[5782] = 14'b0000000_0000000;
		Dplus[5783] = 14'b0000000_0000000;
		Dplus[5784] = 14'b0000000_0000000;
		Dplus[5785] = 14'b0000000_0000000;
		Dplus[5786] = 14'b0000000_0000000;
		Dplus[5787] = 14'b0000000_0000000;
		Dplus[5788] = 14'b0000000_0000000;
		Dplus[5789] = 14'b0000000_0000000;
		Dplus[5790] = 14'b0000000_0000000;
		Dplus[5791] = 14'b0000000_0000000;
		Dplus[5792] = 14'b0000000_0000000;
		Dplus[5793] = 14'b0000000_0000000;
		Dplus[5794] = 14'b0000000_0000000;
		Dplus[5795] = 14'b0000000_0000000;
		Dplus[5796] = 14'b0000000_0000000;
		Dplus[5797] = 14'b0000000_0000000;
		Dplus[5798] = 14'b0000000_0000000;
		Dplus[5799] = 14'b0000000_0000000;
		Dplus[5800] = 14'b0000000_0000000;
		Dplus[5801] = 14'b0000000_0000000;
		Dplus[5802] = 14'b0000000_0000000;
		Dplus[5803] = 14'b0000000_0000000;
		Dplus[5804] = 14'b0000000_0000000;
		Dplus[5805] = 14'b0000000_0000000;
		Dplus[5806] = 14'b0000000_0000000;
		Dplus[5807] = 14'b0000000_0000000;
		Dplus[5808] = 14'b0000000_0000000;
		Dplus[5809] = 14'b0000000_0000000;
		Dplus[5810] = 14'b0000000_0000000;
		Dplus[5811] = 14'b0000000_0000000;
		Dplus[5812] = 14'b0000000_0000000;
		Dplus[5813] = 14'b0000000_0000000;
		Dplus[5814] = 14'b0000000_0000000;
		Dplus[5815] = 14'b0000000_0000000;
		Dplus[5816] = 14'b0000000_0000000;
		Dplus[5817] = 14'b0000000_0000000;
		Dplus[5818] = 14'b0000000_0000000;
		Dplus[5819] = 14'b0000000_0000000;
		Dplus[5820] = 14'b0000000_0000000;
		Dplus[5821] = 14'b0000000_0000000;
		Dplus[5822] = 14'b0000000_0000000;
		Dplus[5823] = 14'b0000000_0000000;
		Dplus[5824] = 14'b0000000_0000000;
		Dplus[5825] = 14'b0000000_0000000;
		Dplus[5826] = 14'b0000000_0000000;
		Dplus[5827] = 14'b0000000_0000000;
		Dplus[5828] = 14'b0000000_0000000;
		Dplus[5829] = 14'b0000000_0000000;
		Dplus[5830] = 14'b0000000_0000000;
		Dplus[5831] = 14'b0000000_0000000;
		Dplus[5832] = 14'b0000000_0000000;
		Dplus[5833] = 14'b0000000_0000000;
		Dplus[5834] = 14'b0000000_0000000;
		Dplus[5835] = 14'b0000000_0000000;
		Dplus[5836] = 14'b0000000_0000000;
		Dplus[5837] = 14'b0000000_0000000;
		Dplus[5838] = 14'b0000000_0000000;
		Dplus[5839] = 14'b0000000_0000000;
		Dplus[5840] = 14'b0000000_0000000;
		Dplus[5841] = 14'b0000000_0000000;
		Dplus[5842] = 14'b0000000_0000000;
		Dplus[5843] = 14'b0000000_0000000;
		Dplus[5844] = 14'b0000000_0000000;
		Dplus[5845] = 14'b0000000_0000000;
		Dplus[5846] = 14'b0000000_0000000;
		Dplus[5847] = 14'b0000000_0000000;
		Dplus[5848] = 14'b0000000_0000000;
		Dplus[5849] = 14'b0000000_0000000;
		Dplus[5850] = 14'b0000000_0000000;
		Dplus[5851] = 14'b0000000_0000000;
		Dplus[5852] = 14'b0000000_0000000;
		Dplus[5853] = 14'b0000000_0000000;
		Dplus[5854] = 14'b0000000_0000000;
		Dplus[5855] = 14'b0000000_0000000;
		Dplus[5856] = 14'b0000000_0000000;
		Dplus[5857] = 14'b0000000_0000000;
		Dplus[5858] = 14'b0000000_0000000;
		Dplus[5859] = 14'b0000000_0000000;
		Dplus[5860] = 14'b0000000_0000000;
		Dplus[5861] = 14'b0000000_0000000;
		Dplus[5862] = 14'b0000000_0000000;
		Dplus[5863] = 14'b0000000_0000000;
		Dplus[5864] = 14'b0000000_0000000;
		Dplus[5865] = 14'b0000000_0000000;
		Dplus[5866] = 14'b0000000_0000000;
		Dplus[5867] = 14'b0000000_0000000;
		Dplus[5868] = 14'b0000000_0000000;
		Dplus[5869] = 14'b0000000_0000000;
		Dplus[5870] = 14'b0000000_0000000;
		Dplus[5871] = 14'b0000000_0000000;
		Dplus[5872] = 14'b0000000_0000000;
		Dplus[5873] = 14'b0000000_0000000;
		Dplus[5874] = 14'b0000000_0000000;
		Dplus[5875] = 14'b0000000_0000000;
		Dplus[5876] = 14'b0000000_0000000;
		Dplus[5877] = 14'b0000000_0000000;
		Dplus[5878] = 14'b0000000_0000000;
		Dplus[5879] = 14'b0000000_0000000;
		Dplus[5880] = 14'b0000000_0000000;
		Dplus[5881] = 14'b0000000_0000000;
		Dplus[5882] = 14'b0000000_0000000;
		Dplus[5883] = 14'b0000000_0000000;
		Dplus[5884] = 14'b0000000_0000000;
		Dplus[5885] = 14'b0000000_0000000;
		Dplus[5886] = 14'b0000000_0000000;
		Dplus[5887] = 14'b0000000_0000000;
		Dplus[5888] = 14'b0000000_0000000;
		Dplus[5889] = 14'b0000000_0000000;
		Dplus[5890] = 14'b0000000_0000000;
		Dplus[5891] = 14'b0000000_0000000;
		Dplus[5892] = 14'b0000000_0000000;
		Dplus[5893] = 14'b0000000_0000000;
		Dplus[5894] = 14'b0000000_0000000;
		Dplus[5895] = 14'b0000000_0000000;
		Dplus[5896] = 14'b0000000_0000000;
		Dplus[5897] = 14'b0000000_0000000;
		Dplus[5898] = 14'b0000000_0000000;
		Dplus[5899] = 14'b0000000_0000000;
		Dplus[5900] = 14'b0000000_0000000;
		Dplus[5901] = 14'b0000000_0000000;
		Dplus[5902] = 14'b0000000_0000000;
		Dplus[5903] = 14'b0000000_0000000;
		Dplus[5904] = 14'b0000000_0000000;
		Dplus[5905] = 14'b0000000_0000000;
		Dplus[5906] = 14'b0000000_0000000;
		Dplus[5907] = 14'b0000000_0000000;
		Dplus[5908] = 14'b0000000_0000000;
		Dplus[5909] = 14'b0000000_0000000;
		Dplus[5910] = 14'b0000000_0000000;
		Dplus[5911] = 14'b0000000_0000000;
		Dplus[5912] = 14'b0000000_0000000;
		Dplus[5913] = 14'b0000000_0000000;
		Dplus[5914] = 14'b0000000_0000000;
		Dplus[5915] = 14'b0000000_0000000;
		Dplus[5916] = 14'b0000000_0000000;
		Dplus[5917] = 14'b0000000_0000000;
		Dplus[5918] = 14'b0000000_0000000;
		Dplus[5919] = 14'b0000000_0000000;
		Dplus[5920] = 14'b0000000_0000000;
		Dplus[5921] = 14'b0000000_0000000;
		Dplus[5922] = 14'b0000000_0000000;
		Dplus[5923] = 14'b0000000_0000000;
		Dplus[5924] = 14'b0000000_0000000;
		Dplus[5925] = 14'b0000000_0000000;
		Dplus[5926] = 14'b0000000_0000000;
		Dplus[5927] = 14'b0000000_0000000;
		Dplus[5928] = 14'b0000000_0000000;
		Dplus[5929] = 14'b0000000_0000000;
		Dplus[5930] = 14'b0000000_0000000;
		Dplus[5931] = 14'b0000000_0000000;
		Dplus[5932] = 14'b0000000_0000000;
		Dplus[5933] = 14'b0000000_0000000;
		Dplus[5934] = 14'b0000000_0000000;
		Dplus[5935] = 14'b0000000_0000000;
		Dplus[5936] = 14'b0000000_0000000;
		Dplus[5937] = 14'b0000000_0000000;
		Dplus[5938] = 14'b0000000_0000000;
		Dplus[5939] = 14'b0000000_0000000;
		Dplus[5940] = 14'b0000000_0000000;
		Dplus[5941] = 14'b0000000_0000000;
		Dplus[5942] = 14'b0000000_0000000;
		Dplus[5943] = 14'b0000000_0000000;
		Dplus[5944] = 14'b0000000_0000000;
		Dplus[5945] = 14'b0000000_0000000;
		Dplus[5946] = 14'b0000000_0000000;
		Dplus[5947] = 14'b0000000_0000000;
		Dplus[5948] = 14'b0000000_0000000;
		Dplus[5949] = 14'b0000000_0000000;
		Dplus[5950] = 14'b0000000_0000000;
		Dplus[5951] = 14'b0000000_0000000;
		Dplus[5952] = 14'b0000000_0000000;
		Dplus[5953] = 14'b0000000_0000000;
		Dplus[5954] = 14'b0000000_0000000;
		Dplus[5955] = 14'b0000000_0000000;
		Dplus[5956] = 14'b0000000_0000000;
		Dplus[5957] = 14'b0000000_0000000;
		Dplus[5958] = 14'b0000000_0000000;
		Dplus[5959] = 14'b0000000_0000000;
		Dplus[5960] = 14'b0000000_0000000;
		Dplus[5961] = 14'b0000000_0000000;
		Dplus[5962] = 14'b0000000_0000000;
		Dplus[5963] = 14'b0000000_0000000;
		Dplus[5964] = 14'b0000000_0000000;
		Dplus[5965] = 14'b0000000_0000000;
		Dplus[5966] = 14'b0000000_0000000;
		Dplus[5967] = 14'b0000000_0000000;
		Dplus[5968] = 14'b0000000_0000000;
		Dplus[5969] = 14'b0000000_0000000;
		Dplus[5970] = 14'b0000000_0000000;
		Dplus[5971] = 14'b0000000_0000000;
		Dplus[5972] = 14'b0000000_0000000;
		Dplus[5973] = 14'b0000000_0000000;
		Dplus[5974] = 14'b0000000_0000000;
		Dplus[5975] = 14'b0000000_0000000;
		Dplus[5976] = 14'b0000000_0000000;
		Dplus[5977] = 14'b0000000_0000000;
		Dplus[5978] = 14'b0000000_0000000;
		Dplus[5979] = 14'b0000000_0000000;
		Dplus[5980] = 14'b0000000_0000000;
		Dplus[5981] = 14'b0000000_0000000;
		Dplus[5982] = 14'b0000000_0000000;
		Dplus[5983] = 14'b0000000_0000000;
		Dplus[5984] = 14'b0000000_0000000;
		Dplus[5985] = 14'b0000000_0000000;
		Dplus[5986] = 14'b0000000_0000000;
		Dplus[5987] = 14'b0000000_0000000;
		Dplus[5988] = 14'b0000000_0000000;
		Dplus[5989] = 14'b0000000_0000000;
		Dplus[5990] = 14'b0000000_0000000;
		Dplus[5991] = 14'b0000000_0000000;
		Dplus[5992] = 14'b0000000_0000000;
		Dplus[5993] = 14'b0000000_0000000;
		Dplus[5994] = 14'b0000000_0000000;
		Dplus[5995] = 14'b0000000_0000000;
		Dplus[5996] = 14'b0000000_0000000;
		Dplus[5997] = 14'b0000000_0000000;
		Dplus[5998] = 14'b0000000_0000000;
		Dplus[5999] = 14'b0000000_0000000;
		Dplus[6000] = 14'b0000000_0000000;
		Dplus[6001] = 14'b0000000_0000000;
		Dplus[6002] = 14'b0000000_0000000;
		Dplus[6003] = 14'b0000000_0000000;
		Dplus[6004] = 14'b0000000_0000000;
		Dplus[6005] = 14'b0000000_0000000;
		Dplus[6006] = 14'b0000000_0000000;
		Dplus[6007] = 14'b0000000_0000000;
		Dplus[6008] = 14'b0000000_0000000;
		Dplus[6009] = 14'b0000000_0000000;
		Dplus[6010] = 14'b0000000_0000000;
		Dplus[6011] = 14'b0000000_0000000;
		Dplus[6012] = 14'b0000000_0000000;
		Dplus[6013] = 14'b0000000_0000000;
		Dplus[6014] = 14'b0000000_0000000;
		Dplus[6015] = 14'b0000000_0000000;
		Dplus[6016] = 14'b0000000_0000000;
		Dplus[6017] = 14'b0000000_0000000;
		Dplus[6018] = 14'b0000000_0000000;
		Dplus[6019] = 14'b0000000_0000000;
		Dplus[6020] = 14'b0000000_0000000;
		Dplus[6021] = 14'b0000000_0000000;
		Dplus[6022] = 14'b0000000_0000000;
		Dplus[6023] = 14'b0000000_0000000;
		Dplus[6024] = 14'b0000000_0000000;
		Dplus[6025] = 14'b0000000_0000000;
		Dplus[6026] = 14'b0000000_0000000;
		Dplus[6027] = 14'b0000000_0000000;
		Dplus[6028] = 14'b0000000_0000000;
		Dplus[6029] = 14'b0000000_0000000;
		Dplus[6030] = 14'b0000000_0000000;
		Dplus[6031] = 14'b0000000_0000000;
		Dplus[6032] = 14'b0000000_0000000;
		Dplus[6033] = 14'b0000000_0000000;
		Dplus[6034] = 14'b0000000_0000000;
		Dplus[6035] = 14'b0000000_0000000;
		Dplus[6036] = 14'b0000000_0000000;
		Dplus[6037] = 14'b0000000_0000000;
		Dplus[6038] = 14'b0000000_0000000;
		Dplus[6039] = 14'b0000000_0000000;
		Dplus[6040] = 14'b0000000_0000000;
		Dplus[6041] = 14'b0000000_0000000;
		Dplus[6042] = 14'b0000000_0000000;
		Dplus[6043] = 14'b0000000_0000000;
		Dplus[6044] = 14'b0000000_0000000;
		Dplus[6045] = 14'b0000000_0000000;
		Dplus[6046] = 14'b0000000_0000000;
		Dplus[6047] = 14'b0000000_0000000;
		Dplus[6048] = 14'b0000000_0000000;
		Dplus[6049] = 14'b0000000_0000000;
		Dplus[6050] = 14'b0000000_0000000;
		Dplus[6051] = 14'b0000000_0000000;
		Dplus[6052] = 14'b0000000_0000000;
		Dplus[6053] = 14'b0000000_0000000;
		Dplus[6054] = 14'b0000000_0000000;
		Dplus[6055] = 14'b0000000_0000000;
		Dplus[6056] = 14'b0000000_0000000;
		Dplus[6057] = 14'b0000000_0000000;
		Dplus[6058] = 14'b0000000_0000000;
		Dplus[6059] = 14'b0000000_0000000;
		Dplus[6060] = 14'b0000000_0000000;
		Dplus[6061] = 14'b0000000_0000000;
		Dplus[6062] = 14'b0000000_0000000;
		Dplus[6063] = 14'b0000000_0000000;
		Dplus[6064] = 14'b0000000_0000000;
		Dplus[6065] = 14'b0000000_0000000;
		Dplus[6066] = 14'b0000000_0000000;
		Dplus[6067] = 14'b0000000_0000000;
		Dplus[6068] = 14'b0000000_0000000;
		Dplus[6069] = 14'b0000000_0000000;
		Dplus[6070] = 14'b0000000_0000000;
		Dplus[6071] = 14'b0000000_0000000;
		Dplus[6072] = 14'b0000000_0000000;
		Dplus[6073] = 14'b0000000_0000000;
		Dplus[6074] = 14'b0000000_0000000;
		Dplus[6075] = 14'b0000000_0000000;
		Dplus[6076] = 14'b0000000_0000000;
		Dplus[6077] = 14'b0000000_0000000;
		Dplus[6078] = 14'b0000000_0000000;
		Dplus[6079] = 14'b0000000_0000000;
		Dplus[6080] = 14'b0000000_0000000;
		Dplus[6081] = 14'b0000000_0000000;
		Dplus[6082] = 14'b0000000_0000000;
		Dplus[6083] = 14'b0000000_0000000;
		Dplus[6084] = 14'b0000000_0000000;
		Dplus[6085] = 14'b0000000_0000000;
		Dplus[6086] = 14'b0000000_0000000;
		Dplus[6087] = 14'b0000000_0000000;
		Dplus[6088] = 14'b0000000_0000000;
		Dplus[6089] = 14'b0000000_0000000;
		Dplus[6090] = 14'b0000000_0000000;
		Dplus[6091] = 14'b0000000_0000000;
		Dplus[6092] = 14'b0000000_0000000;
		Dplus[6093] = 14'b0000000_0000000;
		Dplus[6094] = 14'b0000000_0000000;
		Dplus[6095] = 14'b0000000_0000000;
		Dplus[6096] = 14'b0000000_0000000;
		Dplus[6097] = 14'b0000000_0000000;
		Dplus[6098] = 14'b0000000_0000000;
		Dplus[6099] = 14'b0000000_0000000;
		Dplus[6100] = 14'b0000000_0000000;
		Dplus[6101] = 14'b0000000_0000000;
		Dplus[6102] = 14'b0000000_0000000;
		Dplus[6103] = 14'b0000000_0000000;
		Dplus[6104] = 14'b0000000_0000000;
		Dplus[6105] = 14'b0000000_0000000;
		Dplus[6106] = 14'b0000000_0000000;
		Dplus[6107] = 14'b0000000_0000000;
		Dplus[6108] = 14'b0000000_0000000;
		Dplus[6109] = 14'b0000000_0000000;
		Dplus[6110] = 14'b0000000_0000000;
		Dplus[6111] = 14'b0000000_0000000;
		Dplus[6112] = 14'b0000000_0000000;
		Dplus[6113] = 14'b0000000_0000000;
		Dplus[6114] = 14'b0000000_0000000;
		Dplus[6115] = 14'b0000000_0000000;
		Dplus[6116] = 14'b0000000_0000000;
		Dplus[6117] = 14'b0000000_0000000;
		Dplus[6118] = 14'b0000000_0000000;
		Dplus[6119] = 14'b0000000_0000000;
		Dplus[6120] = 14'b0000000_0000000;
		Dplus[6121] = 14'b0000000_0000000;
		Dplus[6122] = 14'b0000000_0000000;
		Dplus[6123] = 14'b0000000_0000000;
		Dplus[6124] = 14'b0000000_0000000;
		Dplus[6125] = 14'b0000000_0000000;
		Dplus[6126] = 14'b0000000_0000000;
		Dplus[6127] = 14'b0000000_0000000;
		Dplus[6128] = 14'b0000000_0000000;
		Dplus[6129] = 14'b0000000_0000000;
		Dplus[6130] = 14'b0000000_0000000;
		Dplus[6131] = 14'b0000000_0000000;
		Dplus[6132] = 14'b0000000_0000000;
		Dplus[6133] = 14'b0000000_0000000;
		Dplus[6134] = 14'b0000000_0000000;
		Dplus[6135] = 14'b0000000_0000000;
		Dplus[6136] = 14'b0000000_0000000;
		Dplus[6137] = 14'b0000000_0000000;
		Dplus[6138] = 14'b0000000_0000000;
		Dplus[6139] = 14'b0000000_0000000;
		Dplus[6140] = 14'b0000000_0000000;
		Dplus[6141] = 14'b0000000_0000000;
		Dplus[6142] = 14'b0000000_0000000;
		Dplus[6143] = 14'b0000000_0000000;
		Dplus[6144] = 14'b0000000_0000000;
		Dplus[6145] = 14'b0000000_0000000;
		Dplus[6146] = 14'b0000000_0000000;
		Dplus[6147] = 14'b0000000_0000000;
		Dplus[6148] = 14'b0000000_0000000;
		Dplus[6149] = 14'b0000000_0000000;
		Dplus[6150] = 14'b0000000_0000000;
		Dplus[6151] = 14'b0000000_0000000;
		Dplus[6152] = 14'b0000000_0000000;
		Dplus[6153] = 14'b0000000_0000000;
		Dplus[6154] = 14'b0000000_0000000;
		Dplus[6155] = 14'b0000000_0000000;
		Dplus[6156] = 14'b0000000_0000000;
		Dplus[6157] = 14'b0000000_0000000;
		Dplus[6158] = 14'b0000000_0000000;
		Dplus[6159] = 14'b0000000_0000000;
		Dplus[6160] = 14'b0000000_0000000;
		Dplus[6161] = 14'b0000000_0000000;
		Dplus[6162] = 14'b0000000_0000000;
		Dplus[6163] = 14'b0000000_0000000;
		Dplus[6164] = 14'b0000000_0000000;
		Dplus[6165] = 14'b0000000_0000000;
		Dplus[6166] = 14'b0000000_0000000;
		Dplus[6167] = 14'b0000000_0000000;
		Dplus[6168] = 14'b0000000_0000000;
		Dplus[6169] = 14'b0000000_0000000;
		Dplus[6170] = 14'b0000000_0000000;
		Dplus[6171] = 14'b0000000_0000000;
		Dplus[6172] = 14'b0000000_0000000;
		Dplus[6173] = 14'b0000000_0000000;
		Dplus[6174] = 14'b0000000_0000000;
		Dplus[6175] = 14'b0000000_0000000;
		Dplus[6176] = 14'b0000000_0000000;
		Dplus[6177] = 14'b0000000_0000000;
		Dplus[6178] = 14'b0000000_0000000;
		Dplus[6179] = 14'b0000000_0000000;
		Dplus[6180] = 14'b0000000_0000000;
		Dplus[6181] = 14'b0000000_0000000;
		Dplus[6182] = 14'b0000000_0000000;
		Dplus[6183] = 14'b0000000_0000000;
		Dplus[6184] = 14'b0000000_0000000;
		Dplus[6185] = 14'b0000000_0000000;
		Dplus[6186] = 14'b0000000_0000000;
		Dplus[6187] = 14'b0000000_0000000;
		Dplus[6188] = 14'b0000000_0000000;
		Dplus[6189] = 14'b0000000_0000000;
		Dplus[6190] = 14'b0000000_0000000;
		Dplus[6191] = 14'b0000000_0000000;
		Dplus[6192] = 14'b0000000_0000000;
		Dplus[6193] = 14'b0000000_0000000;
		Dplus[6194] = 14'b0000000_0000000;
		Dplus[6195] = 14'b0000000_0000000;
		Dplus[6196] = 14'b0000000_0000000;
		Dplus[6197] = 14'b0000000_0000000;
		Dplus[6198] = 14'b0000000_0000000;
		Dplus[6199] = 14'b0000000_0000000;
		Dplus[6200] = 14'b0000000_0000000;
		Dplus[6201] = 14'b0000000_0000000;
		Dplus[6202] = 14'b0000000_0000000;
		Dplus[6203] = 14'b0000000_0000000;
		Dplus[6204] = 14'b0000000_0000000;
		Dplus[6205] = 14'b0000000_0000000;
		Dplus[6206] = 14'b0000000_0000000;
		Dplus[6207] = 14'b0000000_0000000;
		Dplus[6208] = 14'b0000000_0000000;
		Dplus[6209] = 14'b0000000_0000000;
		Dplus[6210] = 14'b0000000_0000000;
		Dplus[6211] = 14'b0000000_0000000;
		Dplus[6212] = 14'b0000000_0000000;
		Dplus[6213] = 14'b0000000_0000000;
		Dplus[6214] = 14'b0000000_0000000;
		Dplus[6215] = 14'b0000000_0000000;
		Dplus[6216] = 14'b0000000_0000000;
		Dplus[6217] = 14'b0000000_0000000;
		Dplus[6218] = 14'b0000000_0000000;
		Dplus[6219] = 14'b0000000_0000000;
		Dplus[6220] = 14'b0000000_0000000;
		Dplus[6221] = 14'b0000000_0000000;
		Dplus[6222] = 14'b0000000_0000000;
		Dplus[6223] = 14'b0000000_0000000;
		Dplus[6224] = 14'b0000000_0000000;
		Dplus[6225] = 14'b0000000_0000000;
		Dplus[6226] = 14'b0000000_0000000;
		Dplus[6227] = 14'b0000000_0000000;
		Dplus[6228] = 14'b0000000_0000000;
		Dplus[6229] = 14'b0000000_0000000;
		Dplus[6230] = 14'b0000000_0000000;
		Dplus[6231] = 14'b0000000_0000000;
		Dplus[6232] = 14'b0000000_0000000;
		Dplus[6233] = 14'b0000000_0000000;
		Dplus[6234] = 14'b0000000_0000000;
		Dplus[6235] = 14'b0000000_0000000;
		Dplus[6236] = 14'b0000000_0000000;
		Dplus[6237] = 14'b0000000_0000000;
		Dplus[6238] = 14'b0000000_0000000;
		Dplus[6239] = 14'b0000000_0000000;
		Dplus[6240] = 14'b0000000_0000000;
		Dplus[6241] = 14'b0000000_0000000;
		Dplus[6242] = 14'b0000000_0000000;
		Dplus[6243] = 14'b0000000_0000000;
		Dplus[6244] = 14'b0000000_0000000;
		Dplus[6245] = 14'b0000000_0000000;
		Dplus[6246] = 14'b0000000_0000000;
		Dplus[6247] = 14'b0000000_0000000;
		Dplus[6248] = 14'b0000000_0000000;
		Dplus[6249] = 14'b0000000_0000000;
		Dplus[6250] = 14'b0000000_0000000;
		Dplus[6251] = 14'b0000000_0000000;
		Dplus[6252] = 14'b0000000_0000000;
		Dplus[6253] = 14'b0000000_0000000;
		Dplus[6254] = 14'b0000000_0000000;
		Dplus[6255] = 14'b0000000_0000000;
		Dplus[6256] = 14'b0000000_0000000;
		Dplus[6257] = 14'b0000000_0000000;
		Dplus[6258] = 14'b0000000_0000000;
		Dplus[6259] = 14'b0000000_0000000;
		Dplus[6260] = 14'b0000000_0000000;
		Dplus[6261] = 14'b0000000_0000000;
		Dplus[6262] = 14'b0000000_0000000;
		Dplus[6263] = 14'b0000000_0000000;
		Dplus[6264] = 14'b0000000_0000000;
		Dplus[6265] = 14'b0000000_0000000;
		Dplus[6266] = 14'b0000000_0000000;
		Dplus[6267] = 14'b0000000_0000000;
		Dplus[6268] = 14'b0000000_0000000;
		Dplus[6269] = 14'b0000000_0000000;
		Dplus[6270] = 14'b0000000_0000000;
		Dplus[6271] = 14'b0000000_0000000;
		Dplus[6272] = 14'b0000000_0000000;
		Dplus[6273] = 14'b0000000_0000000;
		Dplus[6274] = 14'b0000000_0000000;
		Dplus[6275] = 14'b0000000_0000000;
		Dplus[6276] = 14'b0000000_0000000;
		Dplus[6277] = 14'b0000000_0000000;
		Dplus[6278] = 14'b0000000_0000000;
		Dplus[6279] = 14'b0000000_0000000;
		Dplus[6280] = 14'b0000000_0000000;
		Dplus[6281] = 14'b0000000_0000000;
		Dplus[6282] = 14'b0000000_0000000;
		Dplus[6283] = 14'b0000000_0000000;
		Dplus[6284] = 14'b0000000_0000000;
		Dplus[6285] = 14'b0000000_0000000;
		Dplus[6286] = 14'b0000000_0000000;
		Dplus[6287] = 14'b0000000_0000000;
		Dplus[6288] = 14'b0000000_0000000;
		Dplus[6289] = 14'b0000000_0000000;
		Dplus[6290] = 14'b0000000_0000000;
		Dplus[6291] = 14'b0000000_0000000;
		Dplus[6292] = 14'b0000000_0000000;
		Dplus[6293] = 14'b0000000_0000000;
		Dplus[6294] = 14'b0000000_0000000;
		Dplus[6295] = 14'b0000000_0000000;
		Dplus[6296] = 14'b0000000_0000000;
		Dplus[6297] = 14'b0000000_0000000;
		Dplus[6298] = 14'b0000000_0000000;
		Dplus[6299] = 14'b0000000_0000000;
		Dplus[6300] = 14'b0000000_0000000;
		Dplus[6301] = 14'b0000000_0000000;
		Dplus[6302] = 14'b0000000_0000000;
		Dplus[6303] = 14'b0000000_0000000;
		Dplus[6304] = 14'b0000000_0000000;
		Dplus[6305] = 14'b0000000_0000000;
		Dplus[6306] = 14'b0000000_0000000;
		Dplus[6307] = 14'b0000000_0000000;
		Dplus[6308] = 14'b0000000_0000000;
		Dplus[6309] = 14'b0000000_0000000;
		Dplus[6310] = 14'b0000000_0000000;
		Dplus[6311] = 14'b0000000_0000000;
		Dplus[6312] = 14'b0000000_0000000;
		Dplus[6313] = 14'b0000000_0000000;
		Dplus[6314] = 14'b0000000_0000000;
		Dplus[6315] = 14'b0000000_0000000;
		Dplus[6316] = 14'b0000000_0000000;
		Dplus[6317] = 14'b0000000_0000000;
		Dplus[6318] = 14'b0000000_0000000;
		Dplus[6319] = 14'b0000000_0000000;
		Dplus[6320] = 14'b0000000_0000000;
		Dplus[6321] = 14'b0000000_0000000;
		Dplus[6322] = 14'b0000000_0000000;
		Dplus[6323] = 14'b0000000_0000000;
		Dplus[6324] = 14'b0000000_0000000;
		Dplus[6325] = 14'b0000000_0000000;
		Dplus[6326] = 14'b0000000_0000000;
		Dplus[6327] = 14'b0000000_0000000;
		Dplus[6328] = 14'b0000000_0000000;
		Dplus[6329] = 14'b0000000_0000000;
		Dplus[6330] = 14'b0000000_0000000;
		Dplus[6331] = 14'b0000000_0000000;
		Dplus[6332] = 14'b0000000_0000000;
		Dplus[6333] = 14'b0000000_0000000;
		Dplus[6334] = 14'b0000000_0000000;
		Dplus[6335] = 14'b0000000_0000000;
		Dplus[6336] = 14'b0000000_0000000;
		Dplus[6337] = 14'b0000000_0000000;
		Dplus[6338] = 14'b0000000_0000000;
		Dplus[6339] = 14'b0000000_0000000;
		Dplus[6340] = 14'b0000000_0000000;
		Dplus[6341] = 14'b0000000_0000000;
		Dplus[6342] = 14'b0000000_0000000;
		Dplus[6343] = 14'b0000000_0000000;
		Dplus[6344] = 14'b0000000_0000000;
		Dplus[6345] = 14'b0000000_0000000;
		Dplus[6346] = 14'b0000000_0000000;
		Dplus[6347] = 14'b0000000_0000000;
		Dplus[6348] = 14'b0000000_0000000;
		Dplus[6349] = 14'b0000000_0000000;
		Dplus[6350] = 14'b0000000_0000000;
		Dplus[6351] = 14'b0000000_0000000;
		Dplus[6352] = 14'b0000000_0000000;
		Dplus[6353] = 14'b0000000_0000000;
		Dplus[6354] = 14'b0000000_0000000;
		Dplus[6355] = 14'b0000000_0000000;
		Dplus[6356] = 14'b0000000_0000000;
		Dplus[6357] = 14'b0000000_0000000;
		Dplus[6358] = 14'b0000000_0000000;
		Dplus[6359] = 14'b0000000_0000000;
		Dplus[6360] = 14'b0000000_0000000;
		Dplus[6361] = 14'b0000000_0000000;
		Dplus[6362] = 14'b0000000_0000000;
		Dplus[6363] = 14'b0000000_0000000;
		Dplus[6364] = 14'b0000000_0000000;
		Dplus[6365] = 14'b0000000_0000000;
		Dplus[6366] = 14'b0000000_0000000;
		Dplus[6367] = 14'b0000000_0000000;
		Dplus[6368] = 14'b0000000_0000000;
		Dplus[6369] = 14'b0000000_0000000;
		Dplus[6370] = 14'b0000000_0000000;
		Dplus[6371] = 14'b0000000_0000000;
		Dplus[6372] = 14'b0000000_0000000;
		Dplus[6373] = 14'b0000000_0000000;
		Dplus[6374] = 14'b0000000_0000000;
		Dplus[6375] = 14'b0000000_0000000;
		Dplus[6376] = 14'b0000000_0000000;
		Dplus[6377] = 14'b0000000_0000000;
		Dplus[6378] = 14'b0000000_0000000;
		Dplus[6379] = 14'b0000000_0000000;
		Dplus[6380] = 14'b0000000_0000000;
		Dplus[6381] = 14'b0000000_0000000;
		Dplus[6382] = 14'b0000000_0000000;
		Dplus[6383] = 14'b0000000_0000000;
		Dplus[6384] = 14'b0000000_0000000;
		Dplus[6385] = 14'b0000000_0000000;
		Dplus[6386] = 14'b0000000_0000000;
		Dplus[6387] = 14'b0000000_0000000;
		Dplus[6388] = 14'b0000000_0000000;
		Dplus[6389] = 14'b0000000_0000000;
		Dplus[6390] = 14'b0000000_0000000;
		Dplus[6391] = 14'b0000000_0000000;
		Dplus[6392] = 14'b0000000_0000000;
		Dplus[6393] = 14'b0000000_0000000;
		Dplus[6394] = 14'b0000000_0000000;
		Dplus[6395] = 14'b0000000_0000000;
		Dplus[6396] = 14'b0000000_0000000;
		Dplus[6397] = 14'b0000000_0000000;
		Dplus[6398] = 14'b0000000_0000000;
		Dplus[6399] = 14'b0000000_0000000;
		Dplus[6400] = 14'b0000000_0000000;
		Dplus[6401] = 14'b0000000_0000000;
		Dplus[6402] = 14'b0000000_0000000;
		Dplus[6403] = 14'b0000000_0000000;
		Dplus[6404] = 14'b0000000_0000000;
		Dplus[6405] = 14'b0000000_0000000;
		Dplus[6406] = 14'b0000000_0000000;
		Dplus[6407] = 14'b0000000_0000000;
		Dplus[6408] = 14'b0000000_0000000;
		Dplus[6409] = 14'b0000000_0000000;
		Dplus[6410] = 14'b0000000_0000000;
		Dplus[6411] = 14'b0000000_0000000;
		Dplus[6412] = 14'b0000000_0000000;
		Dplus[6413] = 14'b0000000_0000000;
		Dplus[6414] = 14'b0000000_0000000;
		Dplus[6415] = 14'b0000000_0000000;
		Dplus[6416] = 14'b0000000_0000000;
		Dplus[6417] = 14'b0000000_0000000;
		Dplus[6418] = 14'b0000000_0000000;
		Dplus[6419] = 14'b0000000_0000000;
		Dplus[6420] = 14'b0000000_0000000;
		Dplus[6421] = 14'b0000000_0000000;
		Dplus[6422] = 14'b0000000_0000000;
		Dplus[6423] = 14'b0000000_0000000;
		Dplus[6424] = 14'b0000000_0000000;
		Dplus[6425] = 14'b0000000_0000000;
		Dplus[6426] = 14'b0000000_0000000;
		Dplus[6427] = 14'b0000000_0000000;
		Dplus[6428] = 14'b0000000_0000000;
		Dplus[6429] = 14'b0000000_0000000;
		Dplus[6430] = 14'b0000000_0000000;
		Dplus[6431] = 14'b0000000_0000000;
		Dplus[6432] = 14'b0000000_0000000;
		Dplus[6433] = 14'b0000000_0000000;
		Dplus[6434] = 14'b0000000_0000000;
		Dplus[6435] = 14'b0000000_0000000;
		Dplus[6436] = 14'b0000000_0000000;
		Dplus[6437] = 14'b0000000_0000000;
		Dplus[6438] = 14'b0000000_0000000;
		Dplus[6439] = 14'b0000000_0000000;
		Dplus[6440] = 14'b0000000_0000000;
		Dplus[6441] = 14'b0000000_0000000;
		Dplus[6442] = 14'b0000000_0000000;
		Dplus[6443] = 14'b0000000_0000000;
		Dplus[6444] = 14'b0000000_0000000;
		Dplus[6445] = 14'b0000000_0000000;
		Dplus[6446] = 14'b0000000_0000000;
		Dplus[6447] = 14'b0000000_0000000;
		Dplus[6448] = 14'b0000000_0000000;
		Dplus[6449] = 14'b0000000_0000000;
		Dplus[6450] = 14'b0000000_0000000;
		Dplus[6451] = 14'b0000000_0000000;
		Dplus[6452] = 14'b0000000_0000000;
		Dplus[6453] = 14'b0000000_0000000;
		Dplus[6454] = 14'b0000000_0000000;
		Dplus[6455] = 14'b0000000_0000000;
		Dplus[6456] = 14'b0000000_0000000;
		Dplus[6457] = 14'b0000000_0000000;
		Dplus[6458] = 14'b0000000_0000000;
		Dplus[6459] = 14'b0000000_0000000;
		Dplus[6460] = 14'b0000000_0000000;
		Dplus[6461] = 14'b0000000_0000000;
		Dplus[6462] = 14'b0000000_0000000;
		Dplus[6463] = 14'b0000000_0000000;
		Dplus[6464] = 14'b0000000_0000000;
		Dplus[6465] = 14'b0000000_0000000;
		Dplus[6466] = 14'b0000000_0000000;
		Dplus[6467] = 14'b0000000_0000000;
		Dplus[6468] = 14'b0000000_0000000;
		Dplus[6469] = 14'b0000000_0000000;
		Dplus[6470] = 14'b0000000_0000000;
		Dplus[6471] = 14'b0000000_0000000;
		Dplus[6472] = 14'b0000000_0000000;
		Dplus[6473] = 14'b0000000_0000000;
		Dplus[6474] = 14'b0000000_0000000;
		Dplus[6475] = 14'b0000000_0000000;
		Dplus[6476] = 14'b0000000_0000000;
		Dplus[6477] = 14'b0000000_0000000;
		Dplus[6478] = 14'b0000000_0000000;
		Dplus[6479] = 14'b0000000_0000000;
		Dplus[6480] = 14'b0000000_0000000;
		Dplus[6481] = 14'b0000000_0000000;
		Dplus[6482] = 14'b0000000_0000000;
		Dplus[6483] = 14'b0000000_0000000;
		Dplus[6484] = 14'b0000000_0000000;
		Dplus[6485] = 14'b0000000_0000000;
		Dplus[6486] = 14'b0000000_0000000;
		Dplus[6487] = 14'b0000000_0000000;
		Dplus[6488] = 14'b0000000_0000000;
		Dplus[6489] = 14'b0000000_0000000;
		Dplus[6490] = 14'b0000000_0000000;
		Dplus[6491] = 14'b0000000_0000000;
		Dplus[6492] = 14'b0000000_0000000;
		Dplus[6493] = 14'b0000000_0000000;
		Dplus[6494] = 14'b0000000_0000000;
		Dplus[6495] = 14'b0000000_0000000;
		Dplus[6496] = 14'b0000000_0000000;
		Dplus[6497] = 14'b0000000_0000000;
		Dplus[6498] = 14'b0000000_0000000;
		Dplus[6499] = 14'b0000000_0000000;
		Dplus[6500] = 14'b0000000_0000000;
		Dplus[6501] = 14'b0000000_0000000;
		Dplus[6502] = 14'b0000000_0000000;
		Dplus[6503] = 14'b0000000_0000000;
		Dplus[6504] = 14'b0000000_0000000;
		Dplus[6505] = 14'b0000000_0000000;
		Dplus[6506] = 14'b0000000_0000000;
		Dplus[6507] = 14'b0000000_0000000;
		Dplus[6508] = 14'b0000000_0000000;
		Dplus[6509] = 14'b0000000_0000000;
		Dplus[6510] = 14'b0000000_0000000;
		Dplus[6511] = 14'b0000000_0000000;
		Dplus[6512] = 14'b0000000_0000000;
		Dplus[6513] = 14'b0000000_0000000;
		Dplus[6514] = 14'b0000000_0000000;
		Dplus[6515] = 14'b0000000_0000000;
		Dplus[6516] = 14'b0000000_0000000;
		Dplus[6517] = 14'b0000000_0000000;
		Dplus[6518] = 14'b0000000_0000000;
		Dplus[6519] = 14'b0000000_0000000;
		Dplus[6520] = 14'b0000000_0000000;
		Dplus[6521] = 14'b0000000_0000000;
		Dplus[6522] = 14'b0000000_0000000;
		Dplus[6523] = 14'b0000000_0000000;
		Dplus[6524] = 14'b0000000_0000000;
		Dplus[6525] = 14'b0000000_0000000;
		Dplus[6526] = 14'b0000000_0000000;
		Dplus[6527] = 14'b0000000_0000000;
		Dplus[6528] = 14'b0000000_0000000;
		Dplus[6529] = 14'b0000000_0000000;
		Dplus[6530] = 14'b0000000_0000000;
		Dplus[6531] = 14'b0000000_0000000;
		Dplus[6532] = 14'b0000000_0000000;
		Dplus[6533] = 14'b0000000_0000000;
		Dplus[6534] = 14'b0000000_0000000;
		Dplus[6535] = 14'b0000000_0000000;
		Dplus[6536] = 14'b0000000_0000000;
		Dplus[6537] = 14'b0000000_0000000;
		Dplus[6538] = 14'b0000000_0000000;
		Dplus[6539] = 14'b0000000_0000000;
		Dplus[6540] = 14'b0000000_0000000;
		Dplus[6541] = 14'b0000000_0000000;
		Dplus[6542] = 14'b0000000_0000000;
		Dplus[6543] = 14'b0000000_0000000;
		Dplus[6544] = 14'b0000000_0000000;
		Dplus[6545] = 14'b0000000_0000000;
		Dplus[6546] = 14'b0000000_0000000;
		Dplus[6547] = 14'b0000000_0000000;
		Dplus[6548] = 14'b0000000_0000000;
		Dplus[6549] = 14'b0000000_0000000;
		Dplus[6550] = 14'b0000000_0000000;
		Dplus[6551] = 14'b0000000_0000000;
		Dplus[6552] = 14'b0000000_0000000;
		Dplus[6553] = 14'b0000000_0000000;
		Dplus[6554] = 14'b0000000_0000000;
		Dplus[6555] = 14'b0000000_0000000;
		Dplus[6556] = 14'b0000000_0000000;
		Dplus[6557] = 14'b0000000_0000000;
		Dplus[6558] = 14'b0000000_0000000;
		Dplus[6559] = 14'b0000000_0000000;
		Dplus[6560] = 14'b0000000_0000000;
		Dplus[6561] = 14'b0000000_0000000;
		Dplus[6562] = 14'b0000000_0000000;
		Dplus[6563] = 14'b0000000_0000000;
		Dplus[6564] = 14'b0000000_0000000;
		Dplus[6565] = 14'b0000000_0000000;
		Dplus[6566] = 14'b0000000_0000000;
		Dplus[6567] = 14'b0000000_0000000;
		Dplus[6568] = 14'b0000000_0000000;
		Dplus[6569] = 14'b0000000_0000000;
		Dplus[6570] = 14'b0000000_0000000;
		Dplus[6571] = 14'b0000000_0000000;
		Dplus[6572] = 14'b0000000_0000000;
		Dplus[6573] = 14'b0000000_0000000;
		Dplus[6574] = 14'b0000000_0000000;
		Dplus[6575] = 14'b0000000_0000000;
		Dplus[6576] = 14'b0000000_0000000;
		Dplus[6577] = 14'b0000000_0000000;
		Dplus[6578] = 14'b0000000_0000000;
		Dplus[6579] = 14'b0000000_0000000;
		Dplus[6580] = 14'b0000000_0000000;
		Dplus[6581] = 14'b0000000_0000000;
		Dplus[6582] = 14'b0000000_0000000;
		Dplus[6583] = 14'b0000000_0000000;
		Dplus[6584] = 14'b0000000_0000000;
		Dplus[6585] = 14'b0000000_0000000;
		Dplus[6586] = 14'b0000000_0000000;
		Dplus[6587] = 14'b0000000_0000000;
		Dplus[6588] = 14'b0000000_0000000;
		Dplus[6589] = 14'b0000000_0000000;
		Dplus[6590] = 14'b0000000_0000000;
		Dplus[6591] = 14'b0000000_0000000;
		Dplus[6592] = 14'b0000000_0000000;
		Dplus[6593] = 14'b0000000_0000000;
		Dplus[6594] = 14'b0000000_0000000;
		Dplus[6595] = 14'b0000000_0000000;
		Dplus[6596] = 14'b0000000_0000000;
		Dplus[6597] = 14'b0000000_0000000;
		Dplus[6598] = 14'b0000000_0000000;
		Dplus[6599] = 14'b0000000_0000000;
		Dplus[6600] = 14'b0000000_0000000;
		Dplus[6601] = 14'b0000000_0000000;
		Dplus[6602] = 14'b0000000_0000000;
		Dplus[6603] = 14'b0000000_0000000;
		Dplus[6604] = 14'b0000000_0000000;
		Dplus[6605] = 14'b0000000_0000000;
		Dplus[6606] = 14'b0000000_0000000;
		Dplus[6607] = 14'b0000000_0000000;
		Dplus[6608] = 14'b0000000_0000000;
		Dplus[6609] = 14'b0000000_0000000;
		Dplus[6610] = 14'b0000000_0000000;
		Dplus[6611] = 14'b0000000_0000000;
		Dplus[6612] = 14'b0000000_0000000;
		Dplus[6613] = 14'b0000000_0000000;
		Dplus[6614] = 14'b0000000_0000000;
		Dplus[6615] = 14'b0000000_0000000;
		Dplus[6616] = 14'b0000000_0000000;
		Dplus[6617] = 14'b0000000_0000000;
		Dplus[6618] = 14'b0000000_0000000;
		Dplus[6619] = 14'b0000000_0000000;
		Dplus[6620] = 14'b0000000_0000000;
		Dplus[6621] = 14'b0000000_0000000;
		Dplus[6622] = 14'b0000000_0000000;
		Dplus[6623] = 14'b0000000_0000000;
		Dplus[6624] = 14'b0000000_0000000;
		Dplus[6625] = 14'b0000000_0000000;
		Dplus[6626] = 14'b0000000_0000000;
		Dplus[6627] = 14'b0000000_0000000;
		Dplus[6628] = 14'b0000000_0000000;
		Dplus[6629] = 14'b0000000_0000000;
		Dplus[6630] = 14'b0000000_0000000;
		Dplus[6631] = 14'b0000000_0000000;
		Dplus[6632] = 14'b0000000_0000000;
		Dplus[6633] = 14'b0000000_0000000;
		Dplus[6634] = 14'b0000000_0000000;
		Dplus[6635] = 14'b0000000_0000000;
		Dplus[6636] = 14'b0000000_0000000;
		Dplus[6637] = 14'b0000000_0000000;
		Dplus[6638] = 14'b0000000_0000000;
		Dplus[6639] = 14'b0000000_0000000;
		Dplus[6640] = 14'b0000000_0000000;
		Dplus[6641] = 14'b0000000_0000000;
		Dplus[6642] = 14'b0000000_0000000;
		Dplus[6643] = 14'b0000000_0000000;
		Dplus[6644] = 14'b0000000_0000000;
		Dplus[6645] = 14'b0000000_0000000;
		Dplus[6646] = 14'b0000000_0000000;
		Dplus[6647] = 14'b0000000_0000000;
		Dplus[6648] = 14'b0000000_0000000;
		Dplus[6649] = 14'b0000000_0000000;
		Dplus[6650] = 14'b0000000_0000000;
		Dplus[6651] = 14'b0000000_0000000;
		Dplus[6652] = 14'b0000000_0000000;
		Dplus[6653] = 14'b0000000_0000000;
		Dplus[6654] = 14'b0000000_0000000;
		Dplus[6655] = 14'b0000000_0000000;
		Dplus[6656] = 14'b0000000_0000000;
		Dplus[6657] = 14'b0000000_0000000;
		Dplus[6658] = 14'b0000000_0000000;
		Dplus[6659] = 14'b0000000_0000000;
		Dplus[6660] = 14'b0000000_0000000;
		Dplus[6661] = 14'b0000000_0000000;
		Dplus[6662] = 14'b0000000_0000000;
		Dplus[6663] = 14'b0000000_0000000;
		Dplus[6664] = 14'b0000000_0000000;
		Dplus[6665] = 14'b0000000_0000000;
		Dplus[6666] = 14'b0000000_0000000;
		Dplus[6667] = 14'b0000000_0000000;
		Dplus[6668] = 14'b0000000_0000000;
		Dplus[6669] = 14'b0000000_0000000;
		Dplus[6670] = 14'b0000000_0000000;
		Dplus[6671] = 14'b0000000_0000000;
		Dplus[6672] = 14'b0000000_0000000;
		Dplus[6673] = 14'b0000000_0000000;
		Dplus[6674] = 14'b0000000_0000000;
		Dplus[6675] = 14'b0000000_0000000;
		Dplus[6676] = 14'b0000000_0000000;
		Dplus[6677] = 14'b0000000_0000000;
		Dplus[6678] = 14'b0000000_0000000;
		Dplus[6679] = 14'b0000000_0000000;
		Dplus[6680] = 14'b0000000_0000000;
		Dplus[6681] = 14'b0000000_0000000;
		Dplus[6682] = 14'b0000000_0000000;
		Dplus[6683] = 14'b0000000_0000000;
		Dplus[6684] = 14'b0000000_0000000;
		Dplus[6685] = 14'b0000000_0000000;
		Dplus[6686] = 14'b0000000_0000000;
		Dplus[6687] = 14'b0000000_0000000;
		Dplus[6688] = 14'b0000000_0000000;
		Dplus[6689] = 14'b0000000_0000000;
		Dplus[6690] = 14'b0000000_0000000;
		Dplus[6691] = 14'b0000000_0000000;
		Dplus[6692] = 14'b0000000_0000000;
		Dplus[6693] = 14'b0000000_0000000;
		Dplus[6694] = 14'b0000000_0000000;
		Dplus[6695] = 14'b0000000_0000000;
		Dplus[6696] = 14'b0000000_0000000;
		Dplus[6697] = 14'b0000000_0000000;
		Dplus[6698] = 14'b0000000_0000000;
		Dplus[6699] = 14'b0000000_0000000;
		Dplus[6700] = 14'b0000000_0000000;
		Dplus[6701] = 14'b0000000_0000000;
		Dplus[6702] = 14'b0000000_0000000;
		Dplus[6703] = 14'b0000000_0000000;
		Dplus[6704] = 14'b0000000_0000000;
		Dplus[6705] = 14'b0000000_0000000;
		Dplus[6706] = 14'b0000000_0000000;
		Dplus[6707] = 14'b0000000_0000000;
		Dplus[6708] = 14'b0000000_0000000;
		Dplus[6709] = 14'b0000000_0000000;
		Dplus[6710] = 14'b0000000_0000000;
		Dplus[6711] = 14'b0000000_0000000;
		Dplus[6712] = 14'b0000000_0000000;
		Dplus[6713] = 14'b0000000_0000000;
		Dplus[6714] = 14'b0000000_0000000;
		Dplus[6715] = 14'b0000000_0000000;
		Dplus[6716] = 14'b0000000_0000000;
		Dplus[6717] = 14'b0000000_0000000;
		Dplus[6718] = 14'b0000000_0000000;
		Dplus[6719] = 14'b0000000_0000000;
		Dplus[6720] = 14'b0000000_0000000;
		Dplus[6721] = 14'b0000000_0000000;
		Dplus[6722] = 14'b0000000_0000000;
		Dplus[6723] = 14'b0000000_0000000;
		Dplus[6724] = 14'b0000000_0000000;
		Dplus[6725] = 14'b0000000_0000000;
		Dplus[6726] = 14'b0000000_0000000;
		Dplus[6727] = 14'b0000000_0000000;
		Dplus[6728] = 14'b0000000_0000000;
		Dplus[6729] = 14'b0000000_0000000;
		Dplus[6730] = 14'b0000000_0000000;
		Dplus[6731] = 14'b0000000_0000000;
		Dplus[6732] = 14'b0000000_0000000;
		Dplus[6733] = 14'b0000000_0000000;
		Dplus[6734] = 14'b0000000_0000000;
		Dplus[6735] = 14'b0000000_0000000;
		Dplus[6736] = 14'b0000000_0000000;
		Dplus[6737] = 14'b0000000_0000000;
		Dplus[6738] = 14'b0000000_0000000;
		Dplus[6739] = 14'b0000000_0000000;
		Dplus[6740] = 14'b0000000_0000000;
		Dplus[6741] = 14'b0000000_0000000;
		Dplus[6742] = 14'b0000000_0000000;
		Dplus[6743] = 14'b0000000_0000000;
		Dplus[6744] = 14'b0000000_0000000;
		Dplus[6745] = 14'b0000000_0000000;
		Dplus[6746] = 14'b0000000_0000000;
		Dplus[6747] = 14'b0000000_0000000;
		Dplus[6748] = 14'b0000000_0000000;
		Dplus[6749] = 14'b0000000_0000000;
		Dplus[6750] = 14'b0000000_0000000;
		Dplus[6751] = 14'b0000000_0000000;
		Dplus[6752] = 14'b0000000_0000000;
		Dplus[6753] = 14'b0000000_0000000;
		Dplus[6754] = 14'b0000000_0000000;
		Dplus[6755] = 14'b0000000_0000000;
		Dplus[6756] = 14'b0000000_0000000;
		Dplus[6757] = 14'b0000000_0000000;
		Dplus[6758] = 14'b0000000_0000000;
		Dplus[6759] = 14'b0000000_0000000;
		Dplus[6760] = 14'b0000000_0000000;
		Dplus[6761] = 14'b0000000_0000000;
		Dplus[6762] = 14'b0000000_0000000;
		Dplus[6763] = 14'b0000000_0000000;
		Dplus[6764] = 14'b0000000_0000000;
		Dplus[6765] = 14'b0000000_0000000;
		Dplus[6766] = 14'b0000000_0000000;
		Dplus[6767] = 14'b0000000_0000000;
		Dplus[6768] = 14'b0000000_0000000;
		Dplus[6769] = 14'b0000000_0000000;
		Dplus[6770] = 14'b0000000_0000000;
		Dplus[6771] = 14'b0000000_0000000;
		Dplus[6772] = 14'b0000000_0000000;
		Dplus[6773] = 14'b0000000_0000000;
		Dplus[6774] = 14'b0000000_0000000;
		Dplus[6775] = 14'b0000000_0000000;
		Dplus[6776] = 14'b0000000_0000000;
		Dplus[6777] = 14'b0000000_0000000;
		Dplus[6778] = 14'b0000000_0000000;
		Dplus[6779] = 14'b0000000_0000000;
		Dplus[6780] = 14'b0000000_0000000;
		Dplus[6781] = 14'b0000000_0000000;
		Dplus[6782] = 14'b0000000_0000000;
		Dplus[6783] = 14'b0000000_0000000;
		Dplus[6784] = 14'b0000000_0000000;
		Dplus[6785] = 14'b0000000_0000000;
		Dplus[6786] = 14'b0000000_0000000;
		Dplus[6787] = 14'b0000000_0000000;
		Dplus[6788] = 14'b0000000_0000000;
		Dplus[6789] = 14'b0000000_0000000;
		Dplus[6790] = 14'b0000000_0000000;
		Dplus[6791] = 14'b0000000_0000000;
		Dplus[6792] = 14'b0000000_0000000;
		Dplus[6793] = 14'b0000000_0000000;
		Dplus[6794] = 14'b0000000_0000000;
		Dplus[6795] = 14'b0000000_0000000;
		Dplus[6796] = 14'b0000000_0000000;
		Dplus[6797] = 14'b0000000_0000000;
		Dplus[6798] = 14'b0000000_0000000;
		Dplus[6799] = 14'b0000000_0000000;
		Dplus[6800] = 14'b0000000_0000000;
		Dplus[6801] = 14'b0000000_0000000;
		Dplus[6802] = 14'b0000000_0000000;
		Dplus[6803] = 14'b0000000_0000000;
		Dplus[6804] = 14'b0000000_0000000;
		Dplus[6805] = 14'b0000000_0000000;
		Dplus[6806] = 14'b0000000_0000000;
		Dplus[6807] = 14'b0000000_0000000;
		Dplus[6808] = 14'b0000000_0000000;
		Dplus[6809] = 14'b0000000_0000000;
		Dplus[6810] = 14'b0000000_0000000;
		Dplus[6811] = 14'b0000000_0000000;
		Dplus[6812] = 14'b0000000_0000000;
		Dplus[6813] = 14'b0000000_0000000;
		Dplus[6814] = 14'b0000000_0000000;
		Dplus[6815] = 14'b0000000_0000000;
		Dplus[6816] = 14'b0000000_0000000;
		Dplus[6817] = 14'b0000000_0000000;
		Dplus[6818] = 14'b0000000_0000000;
		Dplus[6819] = 14'b0000000_0000000;
		Dplus[6820] = 14'b0000000_0000000;
		Dplus[6821] = 14'b0000000_0000000;
		Dplus[6822] = 14'b0000000_0000000;
		Dplus[6823] = 14'b0000000_0000000;
		Dplus[6824] = 14'b0000000_0000000;
		Dplus[6825] = 14'b0000000_0000000;
		Dplus[6826] = 14'b0000000_0000000;
		Dplus[6827] = 14'b0000000_0000000;
		Dplus[6828] = 14'b0000000_0000000;
		Dplus[6829] = 14'b0000000_0000000;
		Dplus[6830] = 14'b0000000_0000000;
		Dplus[6831] = 14'b0000000_0000000;
		Dplus[6832] = 14'b0000000_0000000;
		Dplus[6833] = 14'b0000000_0000000;
		Dplus[6834] = 14'b0000000_0000000;
		Dplus[6835] = 14'b0000000_0000000;
		Dplus[6836] = 14'b0000000_0000000;
		Dplus[6837] = 14'b0000000_0000000;
		Dplus[6838] = 14'b0000000_0000000;
		Dplus[6839] = 14'b0000000_0000000;
		Dplus[6840] = 14'b0000000_0000000;
		Dplus[6841] = 14'b0000000_0000000;
		Dplus[6842] = 14'b0000000_0000000;
		Dplus[6843] = 14'b0000000_0000000;
		Dplus[6844] = 14'b0000000_0000000;
		Dplus[6845] = 14'b0000000_0000000;
		Dplus[6846] = 14'b0000000_0000000;
		Dplus[6847] = 14'b0000000_0000000;
		Dplus[6848] = 14'b0000000_0000000;
		Dplus[6849] = 14'b0000000_0000000;
		Dplus[6850] = 14'b0000000_0000000;
		Dplus[6851] = 14'b0000000_0000000;
		Dplus[6852] = 14'b0000000_0000000;
		Dplus[6853] = 14'b0000000_0000000;
		Dplus[6854] = 14'b0000000_0000000;
		Dplus[6855] = 14'b0000000_0000000;
		Dplus[6856] = 14'b0000000_0000000;
		Dplus[6857] = 14'b0000000_0000000;
		Dplus[6858] = 14'b0000000_0000000;
		Dplus[6859] = 14'b0000000_0000000;
		Dplus[6860] = 14'b0000000_0000000;
		Dplus[6861] = 14'b0000000_0000000;
		Dplus[6862] = 14'b0000000_0000000;
		Dplus[6863] = 14'b0000000_0000000;
		Dplus[6864] = 14'b0000000_0000000;
		Dplus[6865] = 14'b0000000_0000000;
		Dplus[6866] = 14'b0000000_0000000;
		Dplus[6867] = 14'b0000000_0000000;
		Dplus[6868] = 14'b0000000_0000000;
		Dplus[6869] = 14'b0000000_0000000;
		Dplus[6870] = 14'b0000000_0000000;
		Dplus[6871] = 14'b0000000_0000000;
		Dplus[6872] = 14'b0000000_0000000;
		Dplus[6873] = 14'b0000000_0000000;
		Dplus[6874] = 14'b0000000_0000000;
		Dplus[6875] = 14'b0000000_0000000;
		Dplus[6876] = 14'b0000000_0000000;
		Dplus[6877] = 14'b0000000_0000000;
		Dplus[6878] = 14'b0000000_0000000;
		Dplus[6879] = 14'b0000000_0000000;
		Dplus[6880] = 14'b0000000_0000000;
		Dplus[6881] = 14'b0000000_0000000;
		Dplus[6882] = 14'b0000000_0000000;
		Dplus[6883] = 14'b0000000_0000000;
		Dplus[6884] = 14'b0000000_0000000;
		Dplus[6885] = 14'b0000000_0000000;
		Dplus[6886] = 14'b0000000_0000000;
		Dplus[6887] = 14'b0000000_0000000;
		Dplus[6888] = 14'b0000000_0000000;
		Dplus[6889] = 14'b0000000_0000000;
		Dplus[6890] = 14'b0000000_0000000;
		Dplus[6891] = 14'b0000000_0000000;
		Dplus[6892] = 14'b0000000_0000000;
		Dplus[6893] = 14'b0000000_0000000;
		Dplus[6894] = 14'b0000000_0000000;
		Dplus[6895] = 14'b0000000_0000000;
		Dplus[6896] = 14'b0000000_0000000;
		Dplus[6897] = 14'b0000000_0000000;
		Dplus[6898] = 14'b0000000_0000000;
		Dplus[6899] = 14'b0000000_0000000;
		Dplus[6900] = 14'b0000000_0000000;
		Dplus[6901] = 14'b0000000_0000000;
		Dplus[6902] = 14'b0000000_0000000;
		Dplus[6903] = 14'b0000000_0000000;
		Dplus[6904] = 14'b0000000_0000000;
		Dplus[6905] = 14'b0000000_0000000;
		Dplus[6906] = 14'b0000000_0000000;
		Dplus[6907] = 14'b0000000_0000000;
		Dplus[6908] = 14'b0000000_0000000;
		Dplus[6909] = 14'b0000000_0000000;
		Dplus[6910] = 14'b0000000_0000000;
		Dplus[6911] = 14'b0000000_0000000;
		Dplus[6912] = 14'b0000000_0000000;
		Dplus[6913] = 14'b0000000_0000000;
		Dplus[6914] = 14'b0000000_0000000;
		Dplus[6915] = 14'b0000000_0000000;
		Dplus[6916] = 14'b0000000_0000000;
		Dplus[6917] = 14'b0000000_0000000;
		Dplus[6918] = 14'b0000000_0000000;
		Dplus[6919] = 14'b0000000_0000000;
		Dplus[6920] = 14'b0000000_0000000;
		Dplus[6921] = 14'b0000000_0000000;
		Dplus[6922] = 14'b0000000_0000000;
		Dplus[6923] = 14'b0000000_0000000;
		Dplus[6924] = 14'b0000000_0000000;
		Dplus[6925] = 14'b0000000_0000000;
		Dplus[6926] = 14'b0000000_0000000;
		Dplus[6927] = 14'b0000000_0000000;
		Dplus[6928] = 14'b0000000_0000000;
		Dplus[6929] = 14'b0000000_0000000;
		Dplus[6930] = 14'b0000000_0000000;
		Dplus[6931] = 14'b0000000_0000000;
		Dplus[6932] = 14'b0000000_0000000;
		Dplus[6933] = 14'b0000000_0000000;
		Dplus[6934] = 14'b0000000_0000000;
		Dplus[6935] = 14'b0000000_0000000;
		Dplus[6936] = 14'b0000000_0000000;
		Dplus[6937] = 14'b0000000_0000000;
		Dplus[6938] = 14'b0000000_0000000;
		Dplus[6939] = 14'b0000000_0000000;
		Dplus[6940] = 14'b0000000_0000000;
		Dplus[6941] = 14'b0000000_0000000;
		Dplus[6942] = 14'b0000000_0000000;
		Dplus[6943] = 14'b0000000_0000000;
		Dplus[6944] = 14'b0000000_0000000;
		Dplus[6945] = 14'b0000000_0000000;
		Dplus[6946] = 14'b0000000_0000000;
		Dplus[6947] = 14'b0000000_0000000;
		Dplus[6948] = 14'b0000000_0000000;
		Dplus[6949] = 14'b0000000_0000000;
		Dplus[6950] = 14'b0000000_0000000;
		Dplus[6951] = 14'b0000000_0000000;
		Dplus[6952] = 14'b0000000_0000000;
		Dplus[6953] = 14'b0000000_0000000;
		Dplus[6954] = 14'b0000000_0000000;
		Dplus[6955] = 14'b0000000_0000000;
		Dplus[6956] = 14'b0000000_0000000;
		Dplus[6957] = 14'b0000000_0000000;
		Dplus[6958] = 14'b0000000_0000000;
		Dplus[6959] = 14'b0000000_0000000;
		Dplus[6960] = 14'b0000000_0000000;
		Dplus[6961] = 14'b0000000_0000000;
		Dplus[6962] = 14'b0000000_0000000;
		Dplus[6963] = 14'b0000000_0000000;
		Dplus[6964] = 14'b0000000_0000000;
		Dplus[6965] = 14'b0000000_0000000;
		Dplus[6966] = 14'b0000000_0000000;
		Dplus[6967] = 14'b0000000_0000000;
		Dplus[6968] = 14'b0000000_0000000;
		Dplus[6969] = 14'b0000000_0000000;
		Dplus[6970] = 14'b0000000_0000000;
		Dplus[6971] = 14'b0000000_0000000;
		Dplus[6972] = 14'b0000000_0000000;
		Dplus[6973] = 14'b0000000_0000000;
		Dplus[6974] = 14'b0000000_0000000;
		Dplus[6975] = 14'b0000000_0000000;
		Dplus[6976] = 14'b0000000_0000000;
		Dplus[6977] = 14'b0000000_0000000;
		Dplus[6978] = 14'b0000000_0000000;
		Dplus[6979] = 14'b0000000_0000000;
		Dplus[6980] = 14'b0000000_0000000;
		Dplus[6981] = 14'b0000000_0000000;
		Dplus[6982] = 14'b0000000_0000000;
		Dplus[6983] = 14'b0000000_0000000;
		Dplus[6984] = 14'b0000000_0000000;
		Dplus[6985] = 14'b0000000_0000000;
		Dplus[6986] = 14'b0000000_0000000;
		Dplus[6987] = 14'b0000000_0000000;
		Dplus[6988] = 14'b0000000_0000000;
		Dplus[6989] = 14'b0000000_0000000;
		Dplus[6990] = 14'b0000000_0000000;
		Dplus[6991] = 14'b0000000_0000000;
		Dplus[6992] = 14'b0000000_0000000;
		Dplus[6993] = 14'b0000000_0000000;
		Dplus[6994] = 14'b0000000_0000000;
		Dplus[6995] = 14'b0000000_0000000;
		Dplus[6996] = 14'b0000000_0000000;
		Dplus[6997] = 14'b0000000_0000000;
		Dplus[6998] = 14'b0000000_0000000;
		Dplus[6999] = 14'b0000000_0000000;
		Dplus[7000] = 14'b0000000_0000000;
		Dplus[7001] = 14'b0000000_0000000;
		Dplus[7002] = 14'b0000000_0000000;
		Dplus[7003] = 14'b0000000_0000000;
		Dplus[7004] = 14'b0000000_0000000;
		Dplus[7005] = 14'b0000000_0000000;
		Dplus[7006] = 14'b0000000_0000000;
		Dplus[7007] = 14'b0000000_0000000;
		Dplus[7008] = 14'b0000000_0000000;
		Dplus[7009] = 14'b0000000_0000000;
		Dplus[7010] = 14'b0000000_0000000;
		Dplus[7011] = 14'b0000000_0000000;
		Dplus[7012] = 14'b0000000_0000000;
		Dplus[7013] = 14'b0000000_0000000;
		Dplus[7014] = 14'b0000000_0000000;
		Dplus[7015] = 14'b0000000_0000000;
		Dplus[7016] = 14'b0000000_0000000;
		Dplus[7017] = 14'b0000000_0000000;
		Dplus[7018] = 14'b0000000_0000000;
		Dplus[7019] = 14'b0000000_0000000;
		Dplus[7020] = 14'b0000000_0000000;
		Dplus[7021] = 14'b0000000_0000000;
		Dplus[7022] = 14'b0000000_0000000;
		Dplus[7023] = 14'b0000000_0000000;
		Dplus[7024] = 14'b0000000_0000000;
		Dplus[7025] = 14'b0000000_0000000;
		Dplus[7026] = 14'b0000000_0000000;
		Dplus[7027] = 14'b0000000_0000000;
		Dplus[7028] = 14'b0000000_0000000;
		Dplus[7029] = 14'b0000000_0000000;
		Dplus[7030] = 14'b0000000_0000000;
		Dplus[7031] = 14'b0000000_0000000;
		Dplus[7032] = 14'b0000000_0000000;
		Dplus[7033] = 14'b0000000_0000000;
		Dplus[7034] = 14'b0000000_0000000;
		Dplus[7035] = 14'b0000000_0000000;
		Dplus[7036] = 14'b0000000_0000000;
		Dplus[7037] = 14'b0000000_0000000;
		Dplus[7038] = 14'b0000000_0000000;
		Dplus[7039] = 14'b0000000_0000000;
		Dplus[7040] = 14'b0000000_0000000;
		Dplus[7041] = 14'b0000000_0000000;
		Dplus[7042] = 14'b0000000_0000000;
		Dplus[7043] = 14'b0000000_0000000;
		Dplus[7044] = 14'b0000000_0000000;
		Dplus[7045] = 14'b0000000_0000000;
		Dplus[7046] = 14'b0000000_0000000;
		Dplus[7047] = 14'b0000000_0000000;
		Dplus[7048] = 14'b0000000_0000000;
		Dplus[7049] = 14'b0000000_0000000;
		Dplus[7050] = 14'b0000000_0000000;
		Dplus[7051] = 14'b0000000_0000000;
		Dplus[7052] = 14'b0000000_0000000;
		Dplus[7053] = 14'b0000000_0000000;
		Dplus[7054] = 14'b0000000_0000000;
		Dplus[7055] = 14'b0000000_0000000;
		Dplus[7056] = 14'b0000000_0000000;
		Dplus[7057] = 14'b0000000_0000000;
		Dplus[7058] = 14'b0000000_0000000;
		Dplus[7059] = 14'b0000000_0000000;
		Dplus[7060] = 14'b0000000_0000000;
		Dplus[7061] = 14'b0000000_0000000;
		Dplus[7062] = 14'b0000000_0000000;
		Dplus[7063] = 14'b0000000_0000000;
		Dplus[7064] = 14'b0000000_0000000;
		Dplus[7065] = 14'b0000000_0000000;
		Dplus[7066] = 14'b0000000_0000000;
		Dplus[7067] = 14'b0000000_0000000;
		Dplus[7068] = 14'b0000000_0000000;
		Dplus[7069] = 14'b0000000_0000000;
		Dplus[7070] = 14'b0000000_0000000;
		Dplus[7071] = 14'b0000000_0000000;
		Dplus[7072] = 14'b0000000_0000000;
		Dplus[7073] = 14'b0000000_0000000;
		Dplus[7074] = 14'b0000000_0000000;
		Dplus[7075] = 14'b0000000_0000000;
		Dplus[7076] = 14'b0000000_0000000;
		Dplus[7077] = 14'b0000000_0000000;
		Dplus[7078] = 14'b0000000_0000000;
		Dplus[7079] = 14'b0000000_0000000;
		Dplus[7080] = 14'b0000000_0000000;
		Dplus[7081] = 14'b0000000_0000000;
		Dplus[7082] = 14'b0000000_0000000;
		Dplus[7083] = 14'b0000000_0000000;
		Dplus[7084] = 14'b0000000_0000000;
		Dplus[7085] = 14'b0000000_0000000;
		Dplus[7086] = 14'b0000000_0000000;
		Dplus[7087] = 14'b0000000_0000000;
		Dplus[7088] = 14'b0000000_0000000;
		Dplus[7089] = 14'b0000000_0000000;
		Dplus[7090] = 14'b0000000_0000000;
		Dplus[7091] = 14'b0000000_0000000;
		Dplus[7092] = 14'b0000000_0000000;
		Dplus[7093] = 14'b0000000_0000000;
		Dplus[7094] = 14'b0000000_0000000;
		Dplus[7095] = 14'b0000000_0000000;
		Dplus[7096] = 14'b0000000_0000000;
		Dplus[7097] = 14'b0000000_0000000;
		Dplus[7098] = 14'b0000000_0000000;
		Dplus[7099] = 14'b0000000_0000000;
		Dplus[7100] = 14'b0000000_0000000;
		Dplus[7101] = 14'b0000000_0000000;
		Dplus[7102] = 14'b0000000_0000000;
		Dplus[7103] = 14'b0000000_0000000;
		Dplus[7104] = 14'b0000000_0000000;
		Dplus[7105] = 14'b0000000_0000000;
		Dplus[7106] = 14'b0000000_0000000;
		Dplus[7107] = 14'b0000000_0000000;
		Dplus[7108] = 14'b0000000_0000000;
		Dplus[7109] = 14'b0000000_0000000;
		Dplus[7110] = 14'b0000000_0000000;
		Dplus[7111] = 14'b0000000_0000000;
		Dplus[7112] = 14'b0000000_0000000;
		Dplus[7113] = 14'b0000000_0000000;
		Dplus[7114] = 14'b0000000_0000000;
		Dplus[7115] = 14'b0000000_0000000;
		Dplus[7116] = 14'b0000000_0000000;
		Dplus[7117] = 14'b0000000_0000000;
		Dplus[7118] = 14'b0000000_0000000;
		Dplus[7119] = 14'b0000000_0000000;
		Dplus[7120] = 14'b0000000_0000000;
		Dplus[7121] = 14'b0000000_0000000;
		Dplus[7122] = 14'b0000000_0000000;
		Dplus[7123] = 14'b0000000_0000000;
		Dplus[7124] = 14'b0000000_0000000;
		Dplus[7125] = 14'b0000000_0000000;
		Dplus[7126] = 14'b0000000_0000000;
		Dplus[7127] = 14'b0000000_0000000;
		Dplus[7128] = 14'b0000000_0000000;
		Dplus[7129] = 14'b0000000_0000000;
		Dplus[7130] = 14'b0000000_0000000;
		Dplus[7131] = 14'b0000000_0000000;
		Dplus[7132] = 14'b0000000_0000000;
		Dplus[7133] = 14'b0000000_0000000;
		Dplus[7134] = 14'b0000000_0000000;
		Dplus[7135] = 14'b0000000_0000000;
		Dplus[7136] = 14'b0000000_0000000;
		Dplus[7137] = 14'b0000000_0000000;
		Dplus[7138] = 14'b0000000_0000000;
		Dplus[7139] = 14'b0000000_0000000;
		Dplus[7140] = 14'b0000000_0000000;
		Dplus[7141] = 14'b0000000_0000000;
		Dplus[7142] = 14'b0000000_0000000;
		Dplus[7143] = 14'b0000000_0000000;
		Dplus[7144] = 14'b0000000_0000000;
		Dplus[7145] = 14'b0000000_0000000;
		Dplus[7146] = 14'b0000000_0000000;
		Dplus[7147] = 14'b0000000_0000000;
		Dplus[7148] = 14'b0000000_0000000;
		Dplus[7149] = 14'b0000000_0000000;
		Dplus[7150] = 14'b0000000_0000000;
		Dplus[7151] = 14'b0000000_0000000;
		Dplus[7152] = 14'b0000000_0000000;
		Dplus[7153] = 14'b0000000_0000000;
		Dplus[7154] = 14'b0000000_0000000;
		Dplus[7155] = 14'b0000000_0000000;
		Dplus[7156] = 14'b0000000_0000000;
		Dplus[7157] = 14'b0000000_0000000;
		Dplus[7158] = 14'b0000000_0000000;
		Dplus[7159] = 14'b0000000_0000000;
		Dplus[7160] = 14'b0000000_0000000;
		Dplus[7161] = 14'b0000000_0000000;
		Dplus[7162] = 14'b0000000_0000000;
		Dplus[7163] = 14'b0000000_0000000;
		Dplus[7164] = 14'b0000000_0000000;
		Dplus[7165] = 14'b0000000_0000000;
		Dplus[7166] = 14'b0000000_0000000;
		Dplus[7167] = 14'b0000000_0000000;
		Dplus[7168] = 14'b0000000_0000000;
		Dplus[7169] = 14'b0000000_0000000;
		Dplus[7170] = 14'b0000000_0000000;
		Dplus[7171] = 14'b0000000_0000000;
		Dplus[7172] = 14'b0000000_0000000;
		Dplus[7173] = 14'b0000000_0000000;
		Dplus[7174] = 14'b0000000_0000000;
		Dplus[7175] = 14'b0000000_0000000;
		Dplus[7176] = 14'b0000000_0000000;
		Dplus[7177] = 14'b0000000_0000000;
		Dplus[7178] = 14'b0000000_0000000;
		Dplus[7179] = 14'b0000000_0000000;
		Dplus[7180] = 14'b0000000_0000000;
		Dplus[7181] = 14'b0000000_0000000;
		Dplus[7182] = 14'b0000000_0000000;
		Dplus[7183] = 14'b0000000_0000000;
		Dplus[7184] = 14'b0000000_0000000;
		Dplus[7185] = 14'b0000000_0000000;
		Dplus[7186] = 14'b0000000_0000000;
		Dplus[7187] = 14'b0000000_0000000;
		Dplus[7188] = 14'b0000000_0000000;
		Dplus[7189] = 14'b0000000_0000000;
		Dplus[7190] = 14'b0000000_0000000;
		Dplus[7191] = 14'b0000000_0000000;
		Dplus[7192] = 14'b0000000_0000000;
		Dplus[7193] = 14'b0000000_0000000;
		Dplus[7194] = 14'b0000000_0000000;
		Dplus[7195] = 14'b0000000_0000000;
		Dplus[7196] = 14'b0000000_0000000;
		Dplus[7197] = 14'b0000000_0000000;
		Dplus[7198] = 14'b0000000_0000000;
		Dplus[7199] = 14'b0000000_0000000;
		Dplus[7200] = 14'b0000000_0000000;
		Dplus[7201] = 14'b0000000_0000000;
		Dplus[7202] = 14'b0000000_0000000;
		Dplus[7203] = 14'b0000000_0000000;
		Dplus[7204] = 14'b0000000_0000000;
		Dplus[7205] = 14'b0000000_0000000;
		Dplus[7206] = 14'b0000000_0000000;
		Dplus[7207] = 14'b0000000_0000000;
		Dplus[7208] = 14'b0000000_0000000;
		Dplus[7209] = 14'b0000000_0000000;
		Dplus[7210] = 14'b0000000_0000000;
		Dplus[7211] = 14'b0000000_0000000;
		Dplus[7212] = 14'b0000000_0000000;
		Dplus[7213] = 14'b0000000_0000000;
		Dplus[7214] = 14'b0000000_0000000;
		Dplus[7215] = 14'b0000000_0000000;
		Dplus[7216] = 14'b0000000_0000000;
		Dplus[7217] = 14'b0000000_0000000;
		Dplus[7218] = 14'b0000000_0000000;
		Dplus[7219] = 14'b0000000_0000000;
		Dplus[7220] = 14'b0000000_0000000;
		Dplus[7221] = 14'b0000000_0000000;
		Dplus[7222] = 14'b0000000_0000000;
		Dplus[7223] = 14'b0000000_0000000;
		Dplus[7224] = 14'b0000000_0000000;
		Dplus[7225] = 14'b0000000_0000000;
		Dplus[7226] = 14'b0000000_0000000;
		Dplus[7227] = 14'b0000000_0000000;
		Dplus[7228] = 14'b0000000_0000000;
		Dplus[7229] = 14'b0000000_0000000;
		Dplus[7230] = 14'b0000000_0000000;
		Dplus[7231] = 14'b0000000_0000000;
		Dplus[7232] = 14'b0000000_0000000;
		Dplus[7233] = 14'b0000000_0000000;
		Dplus[7234] = 14'b0000000_0000000;
		Dplus[7235] = 14'b0000000_0000000;
		Dplus[7236] = 14'b0000000_0000000;
		Dplus[7237] = 14'b0000000_0000000;
		Dplus[7238] = 14'b0000000_0000000;
		Dplus[7239] = 14'b0000000_0000000;
		Dplus[7240] = 14'b0000000_0000000;
		Dplus[7241] = 14'b0000000_0000000;
		Dplus[7242] = 14'b0000000_0000000;
		Dplus[7243] = 14'b0000000_0000000;
		Dplus[7244] = 14'b0000000_0000000;
		Dplus[7245] = 14'b0000000_0000000;
		Dplus[7246] = 14'b0000000_0000000;
		Dplus[7247] = 14'b0000000_0000000;
		Dplus[7248] = 14'b0000000_0000000;
		Dplus[7249] = 14'b0000000_0000000;
		Dplus[7250] = 14'b0000000_0000000;
		Dplus[7251] = 14'b0000000_0000000;
		Dplus[7252] = 14'b0000000_0000000;
		Dplus[7253] = 14'b0000000_0000000;
		Dplus[7254] = 14'b0000000_0000000;
		Dplus[7255] = 14'b0000000_0000000;
		Dplus[7256] = 14'b0000000_0000000;
		Dplus[7257] = 14'b0000000_0000000;
		Dplus[7258] = 14'b0000000_0000000;
		Dplus[7259] = 14'b0000000_0000000;
		Dplus[7260] = 14'b0000000_0000000;
		Dplus[7261] = 14'b0000000_0000000;
		Dplus[7262] = 14'b0000000_0000000;
		Dplus[7263] = 14'b0000000_0000000;
		Dplus[7264] = 14'b0000000_0000000;
		Dplus[7265] = 14'b0000000_0000000;
		Dplus[7266] = 14'b0000000_0000000;
		Dplus[7267] = 14'b0000000_0000000;
		Dplus[7268] = 14'b0000000_0000000;
		Dplus[7269] = 14'b0000000_0000000;
		Dplus[7270] = 14'b0000000_0000000;
		Dplus[7271] = 14'b0000000_0000000;
		Dplus[7272] = 14'b0000000_0000000;
		Dplus[7273] = 14'b0000000_0000000;
		Dplus[7274] = 14'b0000000_0000000;
		Dplus[7275] = 14'b0000000_0000000;
		Dplus[7276] = 14'b0000000_0000000;
		Dplus[7277] = 14'b0000000_0000000;
		Dplus[7278] = 14'b0000000_0000000;
		Dplus[7279] = 14'b0000000_0000000;
		Dplus[7280] = 14'b0000000_0000000;
		Dplus[7281] = 14'b0000000_0000000;
		Dplus[7282] = 14'b0000000_0000000;
		Dplus[7283] = 14'b0000000_0000000;
		Dplus[7284] = 14'b0000000_0000000;
		Dplus[7285] = 14'b0000000_0000000;
		Dplus[7286] = 14'b0000000_0000000;
		Dplus[7287] = 14'b0000000_0000000;
		Dplus[7288] = 14'b0000000_0000000;
		Dplus[7289] = 14'b0000000_0000000;
		Dplus[7290] = 14'b0000000_0000000;
		Dplus[7291] = 14'b0000000_0000000;
		Dplus[7292] = 14'b0000000_0000000;
		Dplus[7293] = 14'b0000000_0000000;
		Dplus[7294] = 14'b0000000_0000000;
		Dplus[7295] = 14'b0000000_0000000;
		Dplus[7296] = 14'b0000000_0000000;
		Dplus[7297] = 14'b0000000_0000000;
		Dplus[7298] = 14'b0000000_0000000;
		Dplus[7299] = 14'b0000000_0000000;
		Dplus[7300] = 14'b0000000_0000000;
		Dplus[7301] = 14'b0000000_0000000;
		Dplus[7302] = 14'b0000000_0000000;
		Dplus[7303] = 14'b0000000_0000000;
		Dplus[7304] = 14'b0000000_0000000;
		Dplus[7305] = 14'b0000000_0000000;
		Dplus[7306] = 14'b0000000_0000000;
		Dplus[7307] = 14'b0000000_0000000;
		Dplus[7308] = 14'b0000000_0000000;
		Dplus[7309] = 14'b0000000_0000000;
		Dplus[7310] = 14'b0000000_0000000;
		Dplus[7311] = 14'b0000000_0000000;
		Dplus[7312] = 14'b0000000_0000000;
		Dplus[7313] = 14'b0000000_0000000;
		Dplus[7314] = 14'b0000000_0000000;
		Dplus[7315] = 14'b0000000_0000000;
		Dplus[7316] = 14'b0000000_0000000;
		Dplus[7317] = 14'b0000000_0000000;
		Dplus[7318] = 14'b0000000_0000000;
		Dplus[7319] = 14'b0000000_0000000;
		Dplus[7320] = 14'b0000000_0000000;
		Dplus[7321] = 14'b0000000_0000000;
		Dplus[7322] = 14'b0000000_0000000;
		Dplus[7323] = 14'b0000000_0000000;
		Dplus[7324] = 14'b0000000_0000000;
		Dplus[7325] = 14'b0000000_0000000;
		Dplus[7326] = 14'b0000000_0000000;
		Dplus[7327] = 14'b0000000_0000000;
		Dplus[7328] = 14'b0000000_0000000;
		Dplus[7329] = 14'b0000000_0000000;
		Dplus[7330] = 14'b0000000_0000000;
		Dplus[7331] = 14'b0000000_0000000;
		Dplus[7332] = 14'b0000000_0000000;
		Dplus[7333] = 14'b0000000_0000000;
		Dplus[7334] = 14'b0000000_0000000;
		Dplus[7335] = 14'b0000000_0000000;
		Dplus[7336] = 14'b0000000_0000000;
		Dplus[7337] = 14'b0000000_0000000;
		Dplus[7338] = 14'b0000000_0000000;
		Dplus[7339] = 14'b0000000_0000000;
		Dplus[7340] = 14'b0000000_0000000;
		Dplus[7341] = 14'b0000000_0000000;
		Dplus[7342] = 14'b0000000_0000000;
		Dplus[7343] = 14'b0000000_0000000;
		Dplus[7344] = 14'b0000000_0000000;
		Dplus[7345] = 14'b0000000_0000000;
		Dplus[7346] = 14'b0000000_0000000;
		Dplus[7347] = 14'b0000000_0000000;
		Dplus[7348] = 14'b0000000_0000000;
		Dplus[7349] = 14'b0000000_0000000;
		Dplus[7350] = 14'b0000000_0000000;
		Dplus[7351] = 14'b0000000_0000000;
		Dplus[7352] = 14'b0000000_0000000;
		Dplus[7353] = 14'b0000000_0000000;
		Dplus[7354] = 14'b0000000_0000000;
		Dplus[7355] = 14'b0000000_0000000;
		Dplus[7356] = 14'b0000000_0000000;
		Dplus[7357] = 14'b0000000_0000000;
		Dplus[7358] = 14'b0000000_0000000;
		Dplus[7359] = 14'b0000000_0000000;
		Dplus[7360] = 14'b0000000_0000000;
		Dplus[7361] = 14'b0000000_0000000;
		Dplus[7362] = 14'b0000000_0000000;
		Dplus[7363] = 14'b0000000_0000000;
		Dplus[7364] = 14'b0000000_0000000;
		Dplus[7365] = 14'b0000000_0000000;
		Dplus[7366] = 14'b0000000_0000000;
		Dplus[7367] = 14'b0000000_0000000;
		Dplus[7368] = 14'b0000000_0000000;
		Dplus[7369] = 14'b0000000_0000000;
		Dplus[7370] = 14'b0000000_0000000;
		Dplus[7371] = 14'b0000000_0000000;
		Dplus[7372] = 14'b0000000_0000000;
		Dplus[7373] = 14'b0000000_0000000;
		Dplus[7374] = 14'b0000000_0000000;
		Dplus[7375] = 14'b0000000_0000000;
		Dplus[7376] = 14'b0000000_0000000;
		Dplus[7377] = 14'b0000000_0000000;
		Dplus[7378] = 14'b0000000_0000000;
		Dplus[7379] = 14'b0000000_0000000;
		Dplus[7380] = 14'b0000000_0000000;
		Dplus[7381] = 14'b0000000_0000000;
		Dplus[7382] = 14'b0000000_0000000;
		Dplus[7383] = 14'b0000000_0000000;
		Dplus[7384] = 14'b0000000_0000000;
		Dplus[7385] = 14'b0000000_0000000;
		Dplus[7386] = 14'b0000000_0000000;
		Dplus[7387] = 14'b0000000_0000000;
		Dplus[7388] = 14'b0000000_0000000;
		Dplus[7389] = 14'b0000000_0000000;
		Dplus[7390] = 14'b0000000_0000000;
		Dplus[7391] = 14'b0000000_0000000;
		Dplus[7392] = 14'b0000000_0000000;
		Dplus[7393] = 14'b0000000_0000000;
		Dplus[7394] = 14'b0000000_0000000;
		Dplus[7395] = 14'b0000000_0000000;
		Dplus[7396] = 14'b0000000_0000000;
		Dplus[7397] = 14'b0000000_0000000;
		Dplus[7398] = 14'b0000000_0000000;
		Dplus[7399] = 14'b0000000_0000000;
		Dplus[7400] = 14'b0000000_0000000;
		Dplus[7401] = 14'b0000000_0000000;
		Dplus[7402] = 14'b0000000_0000000;
		Dplus[7403] = 14'b0000000_0000000;
		Dplus[7404] = 14'b0000000_0000000;
		Dplus[7405] = 14'b0000000_0000000;
		Dplus[7406] = 14'b0000000_0000000;
		Dplus[7407] = 14'b0000000_0000000;
		Dplus[7408] = 14'b0000000_0000000;
		Dplus[7409] = 14'b0000000_0000000;
		Dplus[7410] = 14'b0000000_0000000;
		Dplus[7411] = 14'b0000000_0000000;
		Dplus[7412] = 14'b0000000_0000000;
		Dplus[7413] = 14'b0000000_0000000;
		Dplus[7414] = 14'b0000000_0000000;
		Dplus[7415] = 14'b0000000_0000000;
		Dplus[7416] = 14'b0000000_0000000;
		Dplus[7417] = 14'b0000000_0000000;
		Dplus[7418] = 14'b0000000_0000000;
		Dplus[7419] = 14'b0000000_0000000;
		Dplus[7420] = 14'b0000000_0000000;
		Dplus[7421] = 14'b0000000_0000000;
		Dplus[7422] = 14'b0000000_0000000;
		Dplus[7423] = 14'b0000000_0000000;
		Dplus[7424] = 14'b0000000_0000000;
		Dplus[7425] = 14'b0000000_0000000;
		Dplus[7426] = 14'b0000000_0000000;
		Dplus[7427] = 14'b0000000_0000000;
		Dplus[7428] = 14'b0000000_0000000;
		Dplus[7429] = 14'b0000000_0000000;
		Dplus[7430] = 14'b0000000_0000000;
		Dplus[7431] = 14'b0000000_0000000;
		Dplus[7432] = 14'b0000000_0000000;
		Dplus[7433] = 14'b0000000_0000000;
		Dplus[7434] = 14'b0000000_0000000;
		Dplus[7435] = 14'b0000000_0000000;
		Dplus[7436] = 14'b0000000_0000000;
		Dplus[7437] = 14'b0000000_0000000;
		Dplus[7438] = 14'b0000000_0000000;
		Dplus[7439] = 14'b0000000_0000000;
		Dplus[7440] = 14'b0000000_0000000;
		Dplus[7441] = 14'b0000000_0000000;
		Dplus[7442] = 14'b0000000_0000000;
		Dplus[7443] = 14'b0000000_0000000;
		Dplus[7444] = 14'b0000000_0000000;
		Dplus[7445] = 14'b0000000_0000000;
		Dplus[7446] = 14'b0000000_0000000;
		Dplus[7447] = 14'b0000000_0000000;
		Dplus[7448] = 14'b0000000_0000000;
		Dplus[7449] = 14'b0000000_0000000;
		Dplus[7450] = 14'b0000000_0000000;
		Dplus[7451] = 14'b0000000_0000000;
		Dplus[7452] = 14'b0000000_0000000;
		Dplus[7453] = 14'b0000000_0000000;
		Dplus[7454] = 14'b0000000_0000000;
		Dplus[7455] = 14'b0000000_0000000;
		Dplus[7456] = 14'b0000000_0000000;
		Dplus[7457] = 14'b0000000_0000000;
		Dplus[7458] = 14'b0000000_0000000;
		Dplus[7459] = 14'b0000000_0000000;
		Dplus[7460] = 14'b0000000_0000000;
		Dplus[7461] = 14'b0000000_0000000;
		Dplus[7462] = 14'b0000000_0000000;
		Dplus[7463] = 14'b0000000_0000000;
		Dplus[7464] = 14'b0000000_0000000;
		Dplus[7465] = 14'b0000000_0000000;
		Dplus[7466] = 14'b0000000_0000000;
		Dplus[7467] = 14'b0000000_0000000;
		Dplus[7468] = 14'b0000000_0000000;
		Dplus[7469] = 14'b0000000_0000000;
		Dplus[7470] = 14'b0000000_0000000;
		Dplus[7471] = 14'b0000000_0000000;
		Dplus[7472] = 14'b0000000_0000000;
		Dplus[7473] = 14'b0000000_0000000;
		Dplus[7474] = 14'b0000000_0000000;
		Dplus[7475] = 14'b0000000_0000000;
		Dplus[7476] = 14'b0000000_0000000;
		Dplus[7477] = 14'b0000000_0000000;
		Dplus[7478] = 14'b0000000_0000000;
		Dplus[7479] = 14'b0000000_0000000;
		Dplus[7480] = 14'b0000000_0000000;
		Dplus[7481] = 14'b0000000_0000000;
		Dplus[7482] = 14'b0000000_0000000;
		Dplus[7483] = 14'b0000000_0000000;
		Dplus[7484] = 14'b0000000_0000000;
		Dplus[7485] = 14'b0000000_0000000;
		Dplus[7486] = 14'b0000000_0000000;
		Dplus[7487] = 14'b0000000_0000000;
		Dplus[7488] = 14'b0000000_0000000;
		Dplus[7489] = 14'b0000000_0000000;
		Dplus[7490] = 14'b0000000_0000000;
		Dplus[7491] = 14'b0000000_0000000;
		Dplus[7492] = 14'b0000000_0000000;
		Dplus[7493] = 14'b0000000_0000000;
		Dplus[7494] = 14'b0000000_0000000;
		Dplus[7495] = 14'b0000000_0000000;
		Dplus[7496] = 14'b0000000_0000000;
		Dplus[7497] = 14'b0000000_0000000;
		Dplus[7498] = 14'b0000000_0000000;
		Dplus[7499] = 14'b0000000_0000000;
		Dplus[7500] = 14'b0000000_0000000;
		Dplus[7501] = 14'b0000000_0000000;
		Dplus[7502] = 14'b0000000_0000000;
		Dplus[7503] = 14'b0000000_0000000;
		Dplus[7504] = 14'b0000000_0000000;
		Dplus[7505] = 14'b0000000_0000000;
		Dplus[7506] = 14'b0000000_0000000;
		Dplus[7507] = 14'b0000000_0000000;
		Dplus[7508] = 14'b0000000_0000000;
		Dplus[7509] = 14'b0000000_0000000;
		Dplus[7510] = 14'b0000000_0000000;
		Dplus[7511] = 14'b0000000_0000000;
		Dplus[7512] = 14'b0000000_0000000;
		Dplus[7513] = 14'b0000000_0000000;
		Dplus[7514] = 14'b0000000_0000000;
		Dplus[7515] = 14'b0000000_0000000;
		Dplus[7516] = 14'b0000000_0000000;
		Dplus[7517] = 14'b0000000_0000000;
		Dplus[7518] = 14'b0000000_0000000;
		Dplus[7519] = 14'b0000000_0000000;
		Dplus[7520] = 14'b0000000_0000000;
		Dplus[7521] = 14'b0000000_0000000;
		Dplus[7522] = 14'b0000000_0000000;
		Dplus[7523] = 14'b0000000_0000000;
		Dplus[7524] = 14'b0000000_0000000;
		Dplus[7525] = 14'b0000000_0000000;
		Dplus[7526] = 14'b0000000_0000000;
		Dplus[7527] = 14'b0000000_0000000;
		Dplus[7528] = 14'b0000000_0000000;
		Dplus[7529] = 14'b0000000_0000000;
		Dplus[7530] = 14'b0000000_0000000;
		Dplus[7531] = 14'b0000000_0000000;
		Dplus[7532] = 14'b0000000_0000000;
		Dplus[7533] = 14'b0000000_0000000;
		Dplus[7534] = 14'b0000000_0000000;
		Dplus[7535] = 14'b0000000_0000000;
		Dplus[7536] = 14'b0000000_0000000;
		Dplus[7537] = 14'b0000000_0000000;
		Dplus[7538] = 14'b0000000_0000000;
		Dplus[7539] = 14'b0000000_0000000;
		Dplus[7540] = 14'b0000000_0000000;
		Dplus[7541] = 14'b0000000_0000000;
		Dplus[7542] = 14'b0000000_0000000;
		Dplus[7543] = 14'b0000000_0000000;
		Dplus[7544] = 14'b0000000_0000000;
		Dplus[7545] = 14'b0000000_0000000;
		Dplus[7546] = 14'b0000000_0000000;
		Dplus[7547] = 14'b0000000_0000000;
		Dplus[7548] = 14'b0000000_0000000;
		Dplus[7549] = 14'b0000000_0000000;
		Dplus[7550] = 14'b0000000_0000000;
		Dplus[7551] = 14'b0000000_0000000;
		Dplus[7552] = 14'b0000000_0000000;
		Dplus[7553] = 14'b0000000_0000000;
		Dplus[7554] = 14'b0000000_0000000;
		Dplus[7555] = 14'b0000000_0000000;
		Dplus[7556] = 14'b0000000_0000000;
		Dplus[7557] = 14'b0000000_0000000;
		Dplus[7558] = 14'b0000000_0000000;
		Dplus[7559] = 14'b0000000_0000000;
		Dplus[7560] = 14'b0000000_0000000;
		Dplus[7561] = 14'b0000000_0000000;
		Dplus[7562] = 14'b0000000_0000000;
		Dplus[7563] = 14'b0000000_0000000;
		Dplus[7564] = 14'b0000000_0000000;
		Dplus[7565] = 14'b0000000_0000000;
		Dplus[7566] = 14'b0000000_0000000;
		Dplus[7567] = 14'b0000000_0000000;
		Dplus[7568] = 14'b0000000_0000000;
		Dplus[7569] = 14'b0000000_0000000;
		Dplus[7570] = 14'b0000000_0000000;
		Dplus[7571] = 14'b0000000_0000000;
		Dplus[7572] = 14'b0000000_0000000;
		Dplus[7573] = 14'b0000000_0000000;
		Dplus[7574] = 14'b0000000_0000000;
		Dplus[7575] = 14'b0000000_0000000;
		Dplus[7576] = 14'b0000000_0000000;
		Dplus[7577] = 14'b0000000_0000000;
		Dplus[7578] = 14'b0000000_0000000;
		Dplus[7579] = 14'b0000000_0000000;
		Dplus[7580] = 14'b0000000_0000000;
		Dplus[7581] = 14'b0000000_0000000;
		Dplus[7582] = 14'b0000000_0000000;
		Dplus[7583] = 14'b0000000_0000000;
		Dplus[7584] = 14'b0000000_0000000;
		Dplus[7585] = 14'b0000000_0000000;
		Dplus[7586] = 14'b0000000_0000000;
		Dplus[7587] = 14'b0000000_0000000;
		Dplus[7588] = 14'b0000000_0000000;
		Dplus[7589] = 14'b0000000_0000000;
		Dplus[7590] = 14'b0000000_0000000;
		Dplus[7591] = 14'b0000000_0000000;
		Dplus[7592] = 14'b0000000_0000000;
		Dplus[7593] = 14'b0000000_0000000;
		Dplus[7594] = 14'b0000000_0000000;
		Dplus[7595] = 14'b0000000_0000000;
		Dplus[7596] = 14'b0000000_0000000;
		Dplus[7597] = 14'b0000000_0000000;
		Dplus[7598] = 14'b0000000_0000000;
		Dplus[7599] = 14'b0000000_0000000;
		Dplus[7600] = 14'b0000000_0000000;
		Dplus[7601] = 14'b0000000_0000000;
		Dplus[7602] = 14'b0000000_0000000;
		Dplus[7603] = 14'b0000000_0000000;
		Dplus[7604] = 14'b0000000_0000000;
		Dplus[7605] = 14'b0000000_0000000;
		Dplus[7606] = 14'b0000000_0000000;
		Dplus[7607] = 14'b0000000_0000000;
		Dplus[7608] = 14'b0000000_0000000;
		Dplus[7609] = 14'b0000000_0000000;
		Dplus[7610] = 14'b0000000_0000000;
		Dplus[7611] = 14'b0000000_0000000;
		Dplus[7612] = 14'b0000000_0000000;
		Dplus[7613] = 14'b0000000_0000000;
		Dplus[7614] = 14'b0000000_0000000;
		Dplus[7615] = 14'b0000000_0000000;
		Dplus[7616] = 14'b0000000_0000000;
		Dplus[7617] = 14'b0000000_0000000;
		Dplus[7618] = 14'b0000000_0000000;
		Dplus[7619] = 14'b0000000_0000000;
		Dplus[7620] = 14'b0000000_0000000;
		Dplus[7621] = 14'b0000000_0000000;
		Dplus[7622] = 14'b0000000_0000000;
		Dplus[7623] = 14'b0000000_0000000;
		Dplus[7624] = 14'b0000000_0000000;
		Dplus[7625] = 14'b0000000_0000000;
		Dplus[7626] = 14'b0000000_0000000;
		Dplus[7627] = 14'b0000000_0000000;
		Dplus[7628] = 14'b0000000_0000000;
		Dplus[7629] = 14'b0000000_0000000;
		Dplus[7630] = 14'b0000000_0000000;
		Dplus[7631] = 14'b0000000_0000000;
		Dplus[7632] = 14'b0000000_0000000;
		Dplus[7633] = 14'b0000000_0000000;
		Dplus[7634] = 14'b0000000_0000000;
		Dplus[7635] = 14'b0000000_0000000;
		Dplus[7636] = 14'b0000000_0000000;
		Dplus[7637] = 14'b0000000_0000000;
		Dplus[7638] = 14'b0000000_0000000;
		Dplus[7639] = 14'b0000000_0000000;
		Dplus[7640] = 14'b0000000_0000000;
		Dplus[7641] = 14'b0000000_0000000;
		Dplus[7642] = 14'b0000000_0000000;
		Dplus[7643] = 14'b0000000_0000000;
		Dplus[7644] = 14'b0000000_0000000;
		Dplus[7645] = 14'b0000000_0000000;
		Dplus[7646] = 14'b0000000_0000000;
		Dplus[7647] = 14'b0000000_0000000;
		Dplus[7648] = 14'b0000000_0000000;
		Dplus[7649] = 14'b0000000_0000000;
		Dplus[7650] = 14'b0000000_0000000;
		Dplus[7651] = 14'b0000000_0000000;
		Dplus[7652] = 14'b0000000_0000000;
		Dplus[7653] = 14'b0000000_0000000;
		Dplus[7654] = 14'b0000000_0000000;
		Dplus[7655] = 14'b0000000_0000000;
		Dplus[7656] = 14'b0000000_0000000;
		Dplus[7657] = 14'b0000000_0000000;
		Dplus[7658] = 14'b0000000_0000000;
		Dplus[7659] = 14'b0000000_0000000;
		Dplus[7660] = 14'b0000000_0000000;
		Dplus[7661] = 14'b0000000_0000000;
		Dplus[7662] = 14'b0000000_0000000;
		Dplus[7663] = 14'b0000000_0000000;
		Dplus[7664] = 14'b0000000_0000000;
		Dplus[7665] = 14'b0000000_0000000;
		Dplus[7666] = 14'b0000000_0000000;
		Dplus[7667] = 14'b0000000_0000000;
		Dplus[7668] = 14'b0000000_0000000;
		Dplus[7669] = 14'b0000000_0000000;
		Dplus[7670] = 14'b0000000_0000000;
		Dplus[7671] = 14'b0000000_0000000;
		Dplus[7672] = 14'b0000000_0000000;
		Dplus[7673] = 14'b0000000_0000000;
		Dplus[7674] = 14'b0000000_0000000;
		Dplus[7675] = 14'b0000000_0000000;
		Dplus[7676] = 14'b0000000_0000000;
		Dplus[7677] = 14'b0000000_0000000;
		Dplus[7678] = 14'b0000000_0000000;
		Dplus[7679] = 14'b0000000_0000000;
		Dplus[7680] = 14'b0000000_0000000;
		Dplus[7681] = 14'b0000000_0000000;
		Dplus[7682] = 14'b0000000_0000000;
		Dplus[7683] = 14'b0000000_0000000;
		Dplus[7684] = 14'b0000000_0000000;
		Dplus[7685] = 14'b0000000_0000000;
		Dplus[7686] = 14'b0000000_0000000;
		Dplus[7687] = 14'b0000000_0000000;
		Dplus[7688] = 14'b0000000_0000000;
		Dplus[7689] = 14'b0000000_0000000;
		Dplus[7690] = 14'b0000000_0000000;
		Dplus[7691] = 14'b0000000_0000000;
		Dplus[7692] = 14'b0000000_0000000;
		Dplus[7693] = 14'b0000000_0000000;
		Dplus[7694] = 14'b0000000_0000000;
		Dplus[7695] = 14'b0000000_0000000;
		Dplus[7696] = 14'b0000000_0000000;
		Dplus[7697] = 14'b0000000_0000000;
		Dplus[7698] = 14'b0000000_0000000;
		Dplus[7699] = 14'b0000000_0000000;
		Dplus[7700] = 14'b0000000_0000000;
		Dplus[7701] = 14'b0000000_0000000;
		Dplus[7702] = 14'b0000000_0000000;
		Dplus[7703] = 14'b0000000_0000000;
		Dplus[7704] = 14'b0000000_0000000;
		Dplus[7705] = 14'b0000000_0000000;
		Dplus[7706] = 14'b0000000_0000000;
		Dplus[7707] = 14'b0000000_0000000;
		Dplus[7708] = 14'b0000000_0000000;
		Dplus[7709] = 14'b0000000_0000000;
		Dplus[7710] = 14'b0000000_0000000;
		Dplus[7711] = 14'b0000000_0000000;
		Dplus[7712] = 14'b0000000_0000000;
		Dplus[7713] = 14'b0000000_0000000;
		Dplus[7714] = 14'b0000000_0000000;
		Dplus[7715] = 14'b0000000_0000000;
		Dplus[7716] = 14'b0000000_0000000;
		Dplus[7717] = 14'b0000000_0000000;
		Dplus[7718] = 14'b0000000_0000000;
		Dplus[7719] = 14'b0000000_0000000;
		Dplus[7720] = 14'b0000000_0000000;
		Dplus[7721] = 14'b0000000_0000000;
		Dplus[7722] = 14'b0000000_0000000;
		Dplus[7723] = 14'b0000000_0000000;
		Dplus[7724] = 14'b0000000_0000000;
		Dplus[7725] = 14'b0000000_0000000;
		Dplus[7726] = 14'b0000000_0000000;
		Dplus[7727] = 14'b0000000_0000000;
		Dplus[7728] = 14'b0000000_0000000;
		Dplus[7729] = 14'b0000000_0000000;
		Dplus[7730] = 14'b0000000_0000000;
		Dplus[7731] = 14'b0000000_0000000;
		Dplus[7732] = 14'b0000000_0000000;
		Dplus[7733] = 14'b0000000_0000000;
		Dplus[7734] = 14'b0000000_0000000;
		Dplus[7735] = 14'b0000000_0000000;
		Dplus[7736] = 14'b0000000_0000000;
		Dplus[7737] = 14'b0000000_0000000;
		Dplus[7738] = 14'b0000000_0000000;
		Dplus[7739] = 14'b0000000_0000000;
		Dplus[7740] = 14'b0000000_0000000;
		Dplus[7741] = 14'b0000000_0000000;
		Dplus[7742] = 14'b0000000_0000000;
		Dplus[7743] = 14'b0000000_0000000;
		Dplus[7744] = 14'b0000000_0000000;
		Dplus[7745] = 14'b0000000_0000000;
		Dplus[7746] = 14'b0000000_0000000;
		Dplus[7747] = 14'b0000000_0000000;
		Dplus[7748] = 14'b0000000_0000000;
		Dplus[7749] = 14'b0000000_0000000;
		Dplus[7750] = 14'b0000000_0000000;
		Dplus[7751] = 14'b0000000_0000000;
		Dplus[7752] = 14'b0000000_0000000;
		Dplus[7753] = 14'b0000000_0000000;
		Dplus[7754] = 14'b0000000_0000000;
		Dplus[7755] = 14'b0000000_0000000;
		Dplus[7756] = 14'b0000000_0000000;
		Dplus[7757] = 14'b0000000_0000000;
		Dplus[7758] = 14'b0000000_0000000;
		Dplus[7759] = 14'b0000000_0000000;
		Dplus[7760] = 14'b0000000_0000000;
		Dplus[7761] = 14'b0000000_0000000;
		Dplus[7762] = 14'b0000000_0000000;
		Dplus[7763] = 14'b0000000_0000000;
		Dplus[7764] = 14'b0000000_0000000;
		Dplus[7765] = 14'b0000000_0000000;
		Dplus[7766] = 14'b0000000_0000000;
		Dplus[7767] = 14'b0000000_0000000;
		Dplus[7768] = 14'b0000000_0000000;
		Dplus[7769] = 14'b0000000_0000000;
		Dplus[7770] = 14'b0000000_0000000;
		Dplus[7771] = 14'b0000000_0000000;
		Dplus[7772] = 14'b0000000_0000000;
		Dplus[7773] = 14'b0000000_0000000;
		Dplus[7774] = 14'b0000000_0000000;
		Dplus[7775] = 14'b0000000_0000000;
		Dplus[7776] = 14'b0000000_0000000;
		Dplus[7777] = 14'b0000000_0000000;
		Dplus[7778] = 14'b0000000_0000000;
		Dplus[7779] = 14'b0000000_0000000;
		Dplus[7780] = 14'b0000000_0000000;
		Dplus[7781] = 14'b0000000_0000000;
		Dplus[7782] = 14'b0000000_0000000;
		Dplus[7783] = 14'b0000000_0000000;
		Dplus[7784] = 14'b0000000_0000000;
		Dplus[7785] = 14'b0000000_0000000;
		Dplus[7786] = 14'b0000000_0000000;
		Dplus[7787] = 14'b0000000_0000000;
		Dplus[7788] = 14'b0000000_0000000;
		Dplus[7789] = 14'b0000000_0000000;
		Dplus[7790] = 14'b0000000_0000000;
		Dplus[7791] = 14'b0000000_0000000;
		Dplus[7792] = 14'b0000000_0000000;
		Dplus[7793] = 14'b0000000_0000000;
		Dplus[7794] = 14'b0000000_0000000;
		Dplus[7795] = 14'b0000000_0000000;
		Dplus[7796] = 14'b0000000_0000000;
		Dplus[7797] = 14'b0000000_0000000;
		Dplus[7798] = 14'b0000000_0000000;
		Dplus[7799] = 14'b0000000_0000000;
		Dplus[7800] = 14'b0000000_0000000;
		Dplus[7801] = 14'b0000000_0000000;
		Dplus[7802] = 14'b0000000_0000000;
		Dplus[7803] = 14'b0000000_0000000;
		Dplus[7804] = 14'b0000000_0000000;
		Dplus[7805] = 14'b0000000_0000000;
		Dplus[7806] = 14'b0000000_0000000;
		Dplus[7807] = 14'b0000000_0000000;
		Dplus[7808] = 14'b0000000_0000000;
		Dplus[7809] = 14'b0000000_0000000;
		Dplus[7810] = 14'b0000000_0000000;
		Dplus[7811] = 14'b0000000_0000000;
		Dplus[7812] = 14'b0000000_0000000;
		Dplus[7813] = 14'b0000000_0000000;
		Dplus[7814] = 14'b0000000_0000000;
		Dplus[7815] = 14'b0000000_0000000;
		Dplus[7816] = 14'b0000000_0000000;
		Dplus[7817] = 14'b0000000_0000000;
		Dplus[7818] = 14'b0000000_0000000;
		Dplus[7819] = 14'b0000000_0000000;
		Dplus[7820] = 14'b0000000_0000000;
		Dplus[7821] = 14'b0000000_0000000;
		Dplus[7822] = 14'b0000000_0000000;
		Dplus[7823] = 14'b0000000_0000000;
		Dplus[7824] = 14'b0000000_0000000;
		Dplus[7825] = 14'b0000000_0000000;
		Dplus[7826] = 14'b0000000_0000000;
		Dplus[7827] = 14'b0000000_0000000;
		Dplus[7828] = 14'b0000000_0000000;
		Dplus[7829] = 14'b0000000_0000000;
		Dplus[7830] = 14'b0000000_0000000;
		Dplus[7831] = 14'b0000000_0000000;
		Dplus[7832] = 14'b0000000_0000000;
		Dplus[7833] = 14'b0000000_0000000;
		Dplus[7834] = 14'b0000000_0000000;
		Dplus[7835] = 14'b0000000_0000000;
		Dplus[7836] = 14'b0000000_0000000;
		Dplus[7837] = 14'b0000000_0000000;
		Dplus[7838] = 14'b0000000_0000000;
		Dplus[7839] = 14'b0000000_0000000;
		Dplus[7840] = 14'b0000000_0000000;
		Dplus[7841] = 14'b0000000_0000000;
		Dplus[7842] = 14'b0000000_0000000;
		Dplus[7843] = 14'b0000000_0000000;
		Dplus[7844] = 14'b0000000_0000000;
		Dplus[7845] = 14'b0000000_0000000;
		Dplus[7846] = 14'b0000000_0000000;
		Dplus[7847] = 14'b0000000_0000000;
		Dplus[7848] = 14'b0000000_0000000;
		Dplus[7849] = 14'b0000000_0000000;
		Dplus[7850] = 14'b0000000_0000000;
		Dplus[7851] = 14'b0000000_0000000;
		Dplus[7852] = 14'b0000000_0000000;
		Dplus[7853] = 14'b0000000_0000000;
		Dplus[7854] = 14'b0000000_0000000;
		Dplus[7855] = 14'b0000000_0000000;
		Dplus[7856] = 14'b0000000_0000000;
		Dplus[7857] = 14'b0000000_0000000;
		Dplus[7858] = 14'b0000000_0000000;
		Dplus[7859] = 14'b0000000_0000000;
		Dplus[7860] = 14'b0000000_0000000;
		Dplus[7861] = 14'b0000000_0000000;
		Dplus[7862] = 14'b0000000_0000000;
		Dplus[7863] = 14'b0000000_0000000;
		Dplus[7864] = 14'b0000000_0000000;
		Dplus[7865] = 14'b0000000_0000000;
		Dplus[7866] = 14'b0000000_0000000;
		Dplus[7867] = 14'b0000000_0000000;
		Dplus[7868] = 14'b0000000_0000000;
		Dplus[7869] = 14'b0000000_0000000;
		Dplus[7870] = 14'b0000000_0000000;
		Dplus[7871] = 14'b0000000_0000000;
		Dplus[7872] = 14'b0000000_0000000;
		Dplus[7873] = 14'b0000000_0000000;
		Dplus[7874] = 14'b0000000_0000000;
		Dplus[7875] = 14'b0000000_0000000;
		Dplus[7876] = 14'b0000000_0000000;
		Dplus[7877] = 14'b0000000_0000000;
		Dplus[7878] = 14'b0000000_0000000;
		Dplus[7879] = 14'b0000000_0000000;
		Dplus[7880] = 14'b0000000_0000000;
		Dplus[7881] = 14'b0000000_0000000;
		Dplus[7882] = 14'b0000000_0000000;
		Dplus[7883] = 14'b0000000_0000000;
		Dplus[7884] = 14'b0000000_0000000;
		Dplus[7885] = 14'b0000000_0000000;
		Dplus[7886] = 14'b0000000_0000000;
		Dplus[7887] = 14'b0000000_0000000;
		Dplus[7888] = 14'b0000000_0000000;
		Dplus[7889] = 14'b0000000_0000000;
		Dplus[7890] = 14'b0000000_0000000;
		Dplus[7891] = 14'b0000000_0000000;
		Dplus[7892] = 14'b0000000_0000000;
		Dplus[7893] = 14'b0000000_0000000;
		Dplus[7894] = 14'b0000000_0000000;
		Dplus[7895] = 14'b0000000_0000000;
		Dplus[7896] = 14'b0000000_0000000;
		Dplus[7897] = 14'b0000000_0000000;
		Dplus[7898] = 14'b0000000_0000000;
		Dplus[7899] = 14'b0000000_0000000;
		Dplus[7900] = 14'b0000000_0000000;
		Dplus[7901] = 14'b0000000_0000000;
		Dplus[7902] = 14'b0000000_0000000;
		Dplus[7903] = 14'b0000000_0000000;
		Dplus[7904] = 14'b0000000_0000000;
		Dplus[7905] = 14'b0000000_0000000;
		Dplus[7906] = 14'b0000000_0000000;
		Dplus[7907] = 14'b0000000_0000000;
		Dplus[7908] = 14'b0000000_0000000;
		Dplus[7909] = 14'b0000000_0000000;
		Dplus[7910] = 14'b0000000_0000000;
		Dplus[7911] = 14'b0000000_0000000;
		Dplus[7912] = 14'b0000000_0000000;
		Dplus[7913] = 14'b0000000_0000000;
		Dplus[7914] = 14'b0000000_0000000;
		Dplus[7915] = 14'b0000000_0000000;
		Dplus[7916] = 14'b0000000_0000000;
		Dplus[7917] = 14'b0000000_0000000;
		Dplus[7918] = 14'b0000000_0000000;
		Dplus[7919] = 14'b0000000_0000000;
		Dplus[7920] = 14'b0000000_0000000;
		Dplus[7921] = 14'b0000000_0000000;
		Dplus[7922] = 14'b0000000_0000000;
		Dplus[7923] = 14'b0000000_0000000;
		Dplus[7924] = 14'b0000000_0000000;
		Dplus[7925] = 14'b0000000_0000000;
		Dplus[7926] = 14'b0000000_0000000;
		Dplus[7927] = 14'b0000000_0000000;
		Dplus[7928] = 14'b0000000_0000000;
		Dplus[7929] = 14'b0000000_0000000;
		Dplus[7930] = 14'b0000000_0000000;
		Dplus[7931] = 14'b0000000_0000000;
		Dplus[7932] = 14'b0000000_0000000;
		Dplus[7933] = 14'b0000000_0000000;
		Dplus[7934] = 14'b0000000_0000000;
		Dplus[7935] = 14'b0000000_0000000;
		Dplus[7936] = 14'b0000000_0000000;
		Dplus[7937] = 14'b0000000_0000000;
		Dplus[7938] = 14'b0000000_0000000;
		Dplus[7939] = 14'b0000000_0000000;
		Dplus[7940] = 14'b0000000_0000000;
		Dplus[7941] = 14'b0000000_0000000;
		Dplus[7942] = 14'b0000000_0000000;
		Dplus[7943] = 14'b0000000_0000000;
		Dplus[7944] = 14'b0000000_0000000;
		Dplus[7945] = 14'b0000000_0000000;
		Dplus[7946] = 14'b0000000_0000000;
		Dplus[7947] = 14'b0000000_0000000;
		Dplus[7948] = 14'b0000000_0000000;
		Dplus[7949] = 14'b0000000_0000000;
		Dplus[7950] = 14'b0000000_0000000;
		Dplus[7951] = 14'b0000000_0000000;
		Dplus[7952] = 14'b0000000_0000000;
		Dplus[7953] = 14'b0000000_0000000;
		Dplus[7954] = 14'b0000000_0000000;
		Dplus[7955] = 14'b0000000_0000000;
		Dplus[7956] = 14'b0000000_0000000;
		Dplus[7957] = 14'b0000000_0000000;
		Dplus[7958] = 14'b0000000_0000000;
		Dplus[7959] = 14'b0000000_0000000;
		Dplus[7960] = 14'b0000000_0000000;
		Dplus[7961] = 14'b0000000_0000000;
		Dplus[7962] = 14'b0000000_0000000;
		Dplus[7963] = 14'b0000000_0000000;
		Dplus[7964] = 14'b0000000_0000000;
		Dplus[7965] = 14'b0000000_0000000;
		Dplus[7966] = 14'b0000000_0000000;
		Dplus[7967] = 14'b0000000_0000000;
		Dplus[7968] = 14'b0000000_0000000;
		Dplus[7969] = 14'b0000000_0000000;
		Dplus[7970] = 14'b0000000_0000000;
		Dplus[7971] = 14'b0000000_0000000;
		Dplus[7972] = 14'b0000000_0000000;
		Dplus[7973] = 14'b0000000_0000000;
		Dplus[7974] = 14'b0000000_0000000;
		Dplus[7975] = 14'b0000000_0000000;
		Dplus[7976] = 14'b0000000_0000000;
		Dplus[7977] = 14'b0000000_0000000;
		Dplus[7978] = 14'b0000000_0000000;
		Dplus[7979] = 14'b0000000_0000000;
		Dplus[7980] = 14'b0000000_0000000;
		Dplus[7981] = 14'b0000000_0000000;
		Dplus[7982] = 14'b0000000_0000000;
		Dplus[7983] = 14'b0000000_0000000;
		Dplus[7984] = 14'b0000000_0000000;
		Dplus[7985] = 14'b0000000_0000000;
		Dplus[7986] = 14'b0000000_0000000;
		Dplus[7987] = 14'b0000000_0000000;
		Dplus[7988] = 14'b0000000_0000000;
		Dplus[7989] = 14'b0000000_0000000;
		Dplus[7990] = 14'b0000000_0000000;
		Dplus[7991] = 14'b0000000_0000000;
		Dplus[7992] = 14'b0000000_0000000;
		Dplus[7993] = 14'b0000000_0000000;
		Dplus[7994] = 14'b0000000_0000000;
		Dplus[7995] = 14'b0000000_0000000;
		Dplus[7996] = 14'b0000000_0000000;
		Dplus[7997] = 14'b0000000_0000000;
		Dplus[7998] = 14'b0000000_0000000;
		Dplus[7999] = 14'b0000000_0000000;
		Dplus[8000] = 14'b0000000_0000000;
		Dplus[8001] = 14'b0000000_0000000;
		Dplus[8002] = 14'b0000000_0000000;
		Dplus[8003] = 14'b0000000_0000000;
		Dplus[8004] = 14'b0000000_0000000;
		Dplus[8005] = 14'b0000000_0000000;
		Dplus[8006] = 14'b0000000_0000000;
		Dplus[8007] = 14'b0000000_0000000;
		Dplus[8008] = 14'b0000000_0000000;
		Dplus[8009] = 14'b0000000_0000000;
		Dplus[8010] = 14'b0000000_0000000;
		Dplus[8011] = 14'b0000000_0000000;
		Dplus[8012] = 14'b0000000_0000000;
		Dplus[8013] = 14'b0000000_0000000;
		Dplus[8014] = 14'b0000000_0000000;
		Dplus[8015] = 14'b0000000_0000000;
		Dplus[8016] = 14'b0000000_0000000;
		Dplus[8017] = 14'b0000000_0000000;
		Dplus[8018] = 14'b0000000_0000000;
		Dplus[8019] = 14'b0000000_0000000;
		Dplus[8020] = 14'b0000000_0000000;
		Dplus[8021] = 14'b0000000_0000000;
		Dplus[8022] = 14'b0000000_0000000;
		Dplus[8023] = 14'b0000000_0000000;
		Dplus[8024] = 14'b0000000_0000000;
		Dplus[8025] = 14'b0000000_0000000;
		Dplus[8026] = 14'b0000000_0000000;
		Dplus[8027] = 14'b0000000_0000000;
		Dplus[8028] = 14'b0000000_0000000;
		Dplus[8029] = 14'b0000000_0000000;
		Dplus[8030] = 14'b0000000_0000000;
		Dplus[8031] = 14'b0000000_0000000;
		Dplus[8032] = 14'b0000000_0000000;
		Dplus[8033] = 14'b0000000_0000000;
		Dplus[8034] = 14'b0000000_0000000;
		Dplus[8035] = 14'b0000000_0000000;
		Dplus[8036] = 14'b0000000_0000000;
		Dplus[8037] = 14'b0000000_0000000;
		Dplus[8038] = 14'b0000000_0000000;
		Dplus[8039] = 14'b0000000_0000000;
		Dplus[8040] = 14'b0000000_0000000;
		Dplus[8041] = 14'b0000000_0000000;
		Dplus[8042] = 14'b0000000_0000000;
		Dplus[8043] = 14'b0000000_0000000;
		Dplus[8044] = 14'b0000000_0000000;
		Dplus[8045] = 14'b0000000_0000000;
		Dplus[8046] = 14'b0000000_0000000;
		Dplus[8047] = 14'b0000000_0000000;
		Dplus[8048] = 14'b0000000_0000000;
		Dplus[8049] = 14'b0000000_0000000;
		Dplus[8050] = 14'b0000000_0000000;
		Dplus[8051] = 14'b0000000_0000000;
		Dplus[8052] = 14'b0000000_0000000;
		Dplus[8053] = 14'b0000000_0000000;
		Dplus[8054] = 14'b0000000_0000000;
		Dplus[8055] = 14'b0000000_0000000;
		Dplus[8056] = 14'b0000000_0000000;
		Dplus[8057] = 14'b0000000_0000000;
		Dplus[8058] = 14'b0000000_0000000;
		Dplus[8059] = 14'b0000000_0000000;
		Dplus[8060] = 14'b0000000_0000000;
		Dplus[8061] = 14'b0000000_0000000;
		Dplus[8062] = 14'b0000000_0000000;
		Dplus[8063] = 14'b0000000_0000000;
		Dplus[8064] = 14'b0000000_0000000;
		Dplus[8065] = 14'b0000000_0000000;
		Dplus[8066] = 14'b0000000_0000000;
		Dplus[8067] = 14'b0000000_0000000;
		Dplus[8068] = 14'b0000000_0000000;
		Dplus[8069] = 14'b0000000_0000000;
		Dplus[8070] = 14'b0000000_0000000;
		Dplus[8071] = 14'b0000000_0000000;
		Dplus[8072] = 14'b0000000_0000000;
		Dplus[8073] = 14'b0000000_0000000;
		Dplus[8074] = 14'b0000000_0000000;
		Dplus[8075] = 14'b0000000_0000000;
		Dplus[8076] = 14'b0000000_0000000;
		Dplus[8077] = 14'b0000000_0000000;
		Dplus[8078] = 14'b0000000_0000000;
		Dplus[8079] = 14'b0000000_0000000;
		Dplus[8080] = 14'b0000000_0000000;
		Dplus[8081] = 14'b0000000_0000000;
		Dplus[8082] = 14'b0000000_0000000;
		Dplus[8083] = 14'b0000000_0000000;
		Dplus[8084] = 14'b0000000_0000000;
		Dplus[8085] = 14'b0000000_0000000;
		Dplus[8086] = 14'b0000000_0000000;
		Dplus[8087] = 14'b0000000_0000000;
		Dplus[8088] = 14'b0000000_0000000;
		Dplus[8089] = 14'b0000000_0000000;
		Dplus[8090] = 14'b0000000_0000000;
		Dplus[8091] = 14'b0000000_0000000;
		Dplus[8092] = 14'b0000000_0000000;
		Dplus[8093] = 14'b0000000_0000000;
		Dplus[8094] = 14'b0000000_0000000;
		Dplus[8095] = 14'b0000000_0000000;
		Dplus[8096] = 14'b0000000_0000000;
		Dplus[8097] = 14'b0000000_0000000;
		Dplus[8098] = 14'b0000000_0000000;
		Dplus[8099] = 14'b0000000_0000000;
		Dplus[8100] = 14'b0000000_0000000;
		Dplus[8101] = 14'b0000000_0000000;
		Dplus[8102] = 14'b0000000_0000000;
		Dplus[8103] = 14'b0000000_0000000;
		Dplus[8104] = 14'b0000000_0000000;
		Dplus[8105] = 14'b0000000_0000000;
		Dplus[8106] = 14'b0000000_0000000;
		Dplus[8107] = 14'b0000000_0000000;
		Dplus[8108] = 14'b0000000_0000000;
		Dplus[8109] = 14'b0000000_0000000;
		Dplus[8110] = 14'b0000000_0000000;
		Dplus[8111] = 14'b0000000_0000000;
		Dplus[8112] = 14'b0000000_0000000;
		Dplus[8113] = 14'b0000000_0000000;
		Dplus[8114] = 14'b0000000_0000000;
		Dplus[8115] = 14'b0000000_0000000;
		Dplus[8116] = 14'b0000000_0000000;
		Dplus[8117] = 14'b0000000_0000000;
		Dplus[8118] = 14'b0000000_0000000;
		Dplus[8119] = 14'b0000000_0000000;
		Dplus[8120] = 14'b0000000_0000000;
		Dplus[8121] = 14'b0000000_0000000;
		Dplus[8122] = 14'b0000000_0000000;
		Dplus[8123] = 14'b0000000_0000000;
		Dplus[8124] = 14'b0000000_0000000;
		Dplus[8125] = 14'b0000000_0000000;
		Dplus[8126] = 14'b0000000_0000000;
		Dplus[8127] = 14'b0000000_0000000;
		Dplus[8128] = 14'b0000000_0000000;
		Dplus[8129] = 14'b0000000_0000000;
		Dplus[8130] = 14'b0000000_0000000;
		Dplus[8131] = 14'b0000000_0000000;
		Dplus[8132] = 14'b0000000_0000000;
		Dplus[8133] = 14'b0000000_0000000;
		Dplus[8134] = 14'b0000000_0000000;
		Dplus[8135] = 14'b0000000_0000000;
		Dplus[8136] = 14'b0000000_0000000;
		Dplus[8137] = 14'b0000000_0000000;
		Dplus[8138] = 14'b0000000_0000000;
		Dplus[8139] = 14'b0000000_0000000;
		Dplus[8140] = 14'b0000000_0000000;
		Dplus[8141] = 14'b0000000_0000000;
		Dplus[8142] = 14'b0000000_0000000;
		Dplus[8143] = 14'b0000000_0000000;
		Dplus[8144] = 14'b0000000_0000000;
		Dplus[8145] = 14'b0000000_0000000;
		Dplus[8146] = 14'b0000000_0000000;
		Dplus[8147] = 14'b0000000_0000000;
		Dplus[8148] = 14'b0000000_0000000;
		Dplus[8149] = 14'b0000000_0000000;
		Dplus[8150] = 14'b0000000_0000000;
		Dplus[8151] = 14'b0000000_0000000;
		Dplus[8152] = 14'b0000000_0000000;
		Dplus[8153] = 14'b0000000_0000000;
		Dplus[8154] = 14'b0000000_0000000;
		Dplus[8155] = 14'b0000000_0000000;
		Dplus[8156] = 14'b0000000_0000000;
		Dplus[8157] = 14'b0000000_0000000;
		Dplus[8158] = 14'b0000000_0000000;
		Dplus[8159] = 14'b0000000_0000000;
		Dplus[8160] = 14'b0000000_0000000;
		Dplus[8161] = 14'b0000000_0000000;
		Dplus[8162] = 14'b0000000_0000000;
		Dplus[8163] = 14'b0000000_0000000;
		Dplus[8164] = 14'b0000000_0000000;
		Dplus[8165] = 14'b0000000_0000000;
		Dplus[8166] = 14'b0000000_0000000;
		Dplus[8167] = 14'b0000000_0000000;
		Dplus[8168] = 14'b0000000_0000000;
		Dplus[8169] = 14'b0000000_0000000;
		Dplus[8170] = 14'b0000000_0000000;
		Dplus[8171] = 14'b0000000_0000000;
		Dplus[8172] = 14'b0000000_0000000;
		Dplus[8173] = 14'b0000000_0000000;
		Dplus[8174] = 14'b0000000_0000000;
		Dplus[8175] = 14'b0000000_0000000;
		Dplus[8176] = 14'b0000000_0000000;
		Dplus[8177] = 14'b0000000_0000000;
		Dplus[8178] = 14'b0000000_0000000;
		Dplus[8179] = 14'b0000000_0000000;
		Dplus[8180] = 14'b0000000_0000000;
		Dplus[8181] = 14'b0000000_0000000;
		Dplus[8182] = 14'b0000000_0000000;
		Dplus[8183] = 14'b0000000_0000000;
		Dplus[8184] = 14'b0000000_0000000;
		Dplus[8185] = 14'b0000000_0000000;
		Dplus[8186] = 14'b0000000_0000000;
		Dplus[8187] = 14'b0000000_0000000;
		Dplus[8188] = 14'b0000000_0000000;
		Dplus[8189] = 14'b0000000_0000000;
		Dplus[8190] = 14'b0000000_0000000;
		Dplus[8191] = 14'b0000000_0000000;
end
endmodule
