module Tables();
	reg [9:0] logarithm_table[511:0];
	reg [9:0] Dplus[511:0];
	reg [9:0] Dminus[511:0];
	initial begin
		logarithm_table[1] = 10'b11011_00000;
		logarithm_table[2] = 10'b11100_00000;
		logarithm_table[3] = 10'b11100_10011;
		logarithm_table[4] = 10'b11101_00000;
		logarithm_table[5] = 10'b11101_01010;
		logarithm_table[6] = 10'b11101_10011;
		logarithm_table[7] = 10'b11101_11010;
		logarithm_table[8] = 10'b11110_00000;
		logarithm_table[9] = 10'b11110_00101;
		logarithm_table[10] = 10'b11110_01010;
		logarithm_table[11] = 10'b11110_01111;
		logarithm_table[12] = 10'b11110_10011;
		logarithm_table[13] = 10'b11110_10110;
		logarithm_table[14] = 10'b11110_11010;
		logarithm_table[15] = 10'b11110_11101;
		logarithm_table[16] = 10'b11111_00000;
		logarithm_table[17] = 10'b11111_00011;
		logarithm_table[18] = 10'b11111_00101;
		logarithm_table[19] = 10'b11111_01000;
		logarithm_table[20] = 10'b11111_01010;
		logarithm_table[21] = 10'b11111_01101;
		logarithm_table[22] = 10'b11111_01111;
		logarithm_table[23] = 10'b11111_10001;
		logarithm_table[24] = 10'b11111_10011;
		logarithm_table[25] = 10'b11111_10101;
		logarithm_table[26] = 10'b11111_10110;
		logarithm_table[27] = 10'b11111_11000;
		logarithm_table[28] = 10'b11111_11010;
		logarithm_table[29] = 10'b11111_11011;
		logarithm_table[30] = 10'b11111_11101;
		logarithm_table[31] = 10'b11111_11111;
		logarithm_table[32] = 10'b00000_00000;
		logarithm_table[33] = 10'b00000_00001;
		logarithm_table[34] = 10'b00000_00011;
		logarithm_table[35] = 10'b00000_00100;
		logarithm_table[36] = 10'b00000_00101;
		logarithm_table[37] = 10'b00000_00111;
		logarithm_table[38] = 10'b00000_01000;
		logarithm_table[39] = 10'b00000_01001;
		logarithm_table[40] = 10'b00000_01010;
		logarithm_table[41] = 10'b00000_01011;
		logarithm_table[42] = 10'b00000_01101;
		logarithm_table[43] = 10'b00000_01110;
		logarithm_table[44] = 10'b00000_01111;
		logarithm_table[45] = 10'b00000_10000;
		logarithm_table[46] = 10'b00000_10001;
		logarithm_table[47] = 10'b00000_10010;
		logarithm_table[48] = 10'b00000_10011;
		logarithm_table[49] = 10'b00000_10100;
		logarithm_table[50] = 10'b00000_10101;
		logarithm_table[51] = 10'b00000_10110;
		logarithm_table[52] = 10'b00000_10110;
		logarithm_table[53] = 10'b00000_10111;
		logarithm_table[54] = 10'b00000_11000;
		logarithm_table[55] = 10'b00000_11001;
		logarithm_table[56] = 10'b00000_11010;
		logarithm_table[57] = 10'b00000_11011;
		logarithm_table[58] = 10'b00000_11011;
		logarithm_table[59] = 10'b00000_11100;
		logarithm_table[60] = 10'b00000_11101;
		logarithm_table[61] = 10'b00000_11110;
		logarithm_table[62] = 10'b00000_11111;
		logarithm_table[63] = 10'b00000_11111;
		logarithm_table[64] = 10'b00001_00000;
		logarithm_table[65] = 10'b00001_00001;
		logarithm_table[66] = 10'b00001_00001;
		logarithm_table[67] = 10'b00001_00010;
		logarithm_table[68] = 10'b00001_00011;
		logarithm_table[69] = 10'b00001_00011;
		logarithm_table[70] = 10'b00001_00100;
		logarithm_table[71] = 10'b00001_00101;
		logarithm_table[72] = 10'b00001_00101;
		logarithm_table[73] = 10'b00001_00110;
		logarithm_table[74] = 10'b00001_00111;
		logarithm_table[75] = 10'b00001_00111;
		logarithm_table[76] = 10'b00001_01000;
		logarithm_table[77] = 10'b00001_01001;
		logarithm_table[78] = 10'b00001_01001;
		logarithm_table[79] = 10'b00001_01010;
		logarithm_table[80] = 10'b00001_01010;
		logarithm_table[81] = 10'b00001_01011;
		logarithm_table[82] = 10'b00001_01011;
		logarithm_table[83] = 10'b00001_01100;
		logarithm_table[84] = 10'b00001_01101;
		logarithm_table[85] = 10'b00001_01101;
		logarithm_table[86] = 10'b00001_01110;
		logarithm_table[87] = 10'b00001_01110;
		logarithm_table[88] = 10'b00001_01111;
		logarithm_table[89] = 10'b00001_01111;
		logarithm_table[90] = 10'b00001_10000;
		logarithm_table[91] = 10'b00001_10000;
		logarithm_table[92] = 10'b00001_10001;
		logarithm_table[93] = 10'b00001_10001;
		logarithm_table[94] = 10'b00001_10010;
		logarithm_table[95] = 10'b00001_10010;
		logarithm_table[96] = 10'b00001_10011;
		logarithm_table[97] = 10'b00001_10011;
		logarithm_table[98] = 10'b00001_10100;
		logarithm_table[99] = 10'b00001_10100;
		logarithm_table[100] = 10'b00001_10101;
		logarithm_table[101] = 10'b00001_10101;
		logarithm_table[102] = 10'b00001_10110;
		logarithm_table[103] = 10'b00001_10110;
		logarithm_table[104] = 10'b00001_10110;
		logarithm_table[105] = 10'b00001_10111;
		logarithm_table[106] = 10'b00001_10111;
		logarithm_table[107] = 10'b00001_11000;
		logarithm_table[108] = 10'b00001_11000;
		logarithm_table[109] = 10'b00001_11001;
		logarithm_table[110] = 10'b00001_11001;
		logarithm_table[111] = 10'b00001_11001;
		logarithm_table[112] = 10'b00001_11010;
		logarithm_table[113] = 10'b00001_11010;
		logarithm_table[114] = 10'b00001_11011;
		logarithm_table[115] = 10'b00001_11011;
		logarithm_table[116] = 10'b00001_11011;
		logarithm_table[117] = 10'b00001_11100;
		logarithm_table[118] = 10'b00001_11100;
		logarithm_table[119] = 10'b00001_11101;
		logarithm_table[120] = 10'b00001_11101;
		logarithm_table[121] = 10'b00001_11101;
		logarithm_table[122] = 10'b00001_11110;
		logarithm_table[123] = 10'b00001_11110;
		logarithm_table[124] = 10'b00001_11111;
		logarithm_table[125] = 10'b00001_11111;
		logarithm_table[126] = 10'b00001_11111;
		logarithm_table[127] = 10'b00010_00000;
		logarithm_table[128] = 10'b00010_00000;
		logarithm_table[129] = 10'b00010_00000;
		logarithm_table[130] = 10'b00010_00001;
		logarithm_table[131] = 10'b00010_00001;
		logarithm_table[132] = 10'b00010_00001;
		logarithm_table[133] = 10'b00010_00010;
		logarithm_table[134] = 10'b00010_00010;
		logarithm_table[135] = 10'b00010_00010;
		logarithm_table[136] = 10'b00010_00011;
		logarithm_table[137] = 10'b00010_00011;
		logarithm_table[138] = 10'b00010_00011;
		logarithm_table[139] = 10'b00010_00100;
		logarithm_table[140] = 10'b00010_00100;
		logarithm_table[141] = 10'b00010_00100;
		logarithm_table[142] = 10'b00010_00101;
		logarithm_table[143] = 10'b00010_00101;
		logarithm_table[144] = 10'b00010_00101;
		logarithm_table[145] = 10'b00010_00110;
		logarithm_table[146] = 10'b00010_00110;
		logarithm_table[147] = 10'b00010_00110;
		logarithm_table[148] = 10'b00010_00111;
		logarithm_table[149] = 10'b00010_00111;
		logarithm_table[150] = 10'b00010_00111;
		logarithm_table[151] = 10'b00010_01000;
		logarithm_table[152] = 10'b00010_01000;
		logarithm_table[153] = 10'b00010_01000;
		logarithm_table[154] = 10'b00010_01001;
		logarithm_table[155] = 10'b00010_01001;
		logarithm_table[156] = 10'b00010_01001;
		logarithm_table[157] = 10'b00010_01001;
		logarithm_table[158] = 10'b00010_01010;
		logarithm_table[159] = 10'b00010_01010;
		logarithm_table[160] = 10'b00010_01010;
		logarithm_table[161] = 10'b00010_01011;
		logarithm_table[162] = 10'b00010_01011;
		logarithm_table[163] = 10'b00010_01011;
		logarithm_table[164] = 10'b00010_01011;
		logarithm_table[165] = 10'b00010_01100;
		logarithm_table[166] = 10'b00010_01100;
		logarithm_table[167] = 10'b00010_01100;
		logarithm_table[168] = 10'b00010_01101;
		logarithm_table[169] = 10'b00010_01101;
		logarithm_table[170] = 10'b00010_01101;
		logarithm_table[171] = 10'b00010_01101;
		logarithm_table[172] = 10'b00010_01110;
		logarithm_table[173] = 10'b00010_01110;
		logarithm_table[174] = 10'b00010_01110;
		logarithm_table[175] = 10'b00010_01110;
		logarithm_table[176] = 10'b00010_01111;
		logarithm_table[177] = 10'b00010_01111;
		logarithm_table[178] = 10'b00010_01111;
		logarithm_table[179] = 10'b00010_01111;
		logarithm_table[180] = 10'b00010_10000;
		logarithm_table[181] = 10'b00010_10000;
		logarithm_table[182] = 10'b00010_10000;
		logarithm_table[183] = 10'b00010_10001;
		logarithm_table[184] = 10'b00010_10001;
		logarithm_table[185] = 10'b00010_10001;
		logarithm_table[186] = 10'b00010_10001;
		logarithm_table[187] = 10'b00010_10010;
		logarithm_table[188] = 10'b00010_10010;
		logarithm_table[189] = 10'b00010_10010;
		logarithm_table[190] = 10'b00010_10010;
		logarithm_table[191] = 10'b00010_10010;
		logarithm_table[192] = 10'b00010_10011;
		logarithm_table[193] = 10'b00010_10011;
		logarithm_table[194] = 10'b00010_10011;
		logarithm_table[195] = 10'b00010_10011;
		logarithm_table[196] = 10'b00010_10100;
		logarithm_table[197] = 10'b00010_10100;
		logarithm_table[198] = 10'b00010_10100;
		logarithm_table[199] = 10'b00010_10100;
		logarithm_table[200] = 10'b00010_10101;
		logarithm_table[201] = 10'b00010_10101;
		logarithm_table[202] = 10'b00010_10101;
		logarithm_table[203] = 10'b00010_10101;
		logarithm_table[204] = 10'b00010_10110;
		logarithm_table[205] = 10'b00010_10110;
		logarithm_table[206] = 10'b00010_10110;
		logarithm_table[207] = 10'b00010_10110;
		logarithm_table[208] = 10'b00010_10110;
		logarithm_table[209] = 10'b00010_10111;
		logarithm_table[210] = 10'b00010_10111;
		logarithm_table[211] = 10'b00010_10111;
		logarithm_table[212] = 10'b00010_10111;
		logarithm_table[213] = 10'b00010_11000;
		logarithm_table[214] = 10'b00010_11000;
		logarithm_table[215] = 10'b00010_11000;
		logarithm_table[216] = 10'b00010_11000;
		logarithm_table[217] = 10'b00010_11000;
		logarithm_table[218] = 10'b00010_11001;
		logarithm_table[219] = 10'b00010_11001;
		logarithm_table[220] = 10'b00010_11001;
		logarithm_table[221] = 10'b00010_11001;
		logarithm_table[222] = 10'b00010_11001;
		logarithm_table[223] = 10'b00010_11010;
		logarithm_table[224] = 10'b00010_11010;
		logarithm_table[225] = 10'b00010_11010;
		logarithm_table[226] = 10'b00010_11010;
		logarithm_table[227] = 10'b00010_11010;
		logarithm_table[228] = 10'b00010_11011;
		logarithm_table[229] = 10'b00010_11011;
		logarithm_table[230] = 10'b00010_11011;
		logarithm_table[231] = 10'b00010_11011;
		logarithm_table[232] = 10'b00010_11011;
		logarithm_table[233] = 10'b00010_11100;
		logarithm_table[234] = 10'b00010_11100;
		logarithm_table[235] = 10'b00010_11100;
		logarithm_table[236] = 10'b00010_11100;
		logarithm_table[237] = 10'b00010_11100;
		logarithm_table[238] = 10'b00010_11101;
		logarithm_table[239] = 10'b00010_11101;
		logarithm_table[240] = 10'b00010_11101;
		logarithm_table[241] = 10'b00010_11101;
		logarithm_table[242] = 10'b00010_11101;
		logarithm_table[243] = 10'b00010_11110;
		logarithm_table[244] = 10'b00010_11110;
		logarithm_table[245] = 10'b00010_11110;
		logarithm_table[246] = 10'b00010_11110;
		logarithm_table[247] = 10'b00010_11110;
		logarithm_table[248] = 10'b00010_11111;
		logarithm_table[249] = 10'b00010_11111;
		logarithm_table[250] = 10'b00010_11111;
		logarithm_table[251] = 10'b00010_11111;
		logarithm_table[252] = 10'b00010_11111;
		logarithm_table[253] = 10'b00010_11111;
		logarithm_table[254] = 10'b00011_00000;
		logarithm_table[255] = 10'b00011_00000;
		logarithm_table[256] = 10'b00011_00000;
		logarithm_table[257] = 10'b00011_00000;
		logarithm_table[258] = 10'b00011_00000;
		logarithm_table[259] = 10'b00011_00001;
		logarithm_table[260] = 10'b00011_00001;
		logarithm_table[261] = 10'b00011_00001;
		logarithm_table[262] = 10'b00011_00001;
		logarithm_table[263] = 10'b00011_00001;
		logarithm_table[264] = 10'b00011_00001;
		logarithm_table[265] = 10'b00011_00010;
		logarithm_table[266] = 10'b00011_00010;
		logarithm_table[267] = 10'b00011_00010;
		logarithm_table[268] = 10'b00011_00010;
		logarithm_table[269] = 10'b00011_00010;
		logarithm_table[270] = 10'b00011_00010;
		logarithm_table[271] = 10'b00011_00011;
		logarithm_table[272] = 10'b00011_00011;
		logarithm_table[273] = 10'b00011_00011;
		logarithm_table[274] = 10'b00011_00011;
		logarithm_table[275] = 10'b00011_00011;
		logarithm_table[276] = 10'b00011_00011;
		logarithm_table[277] = 10'b00011_00100;
		logarithm_table[278] = 10'b00011_00100;
		logarithm_table[279] = 10'b00011_00100;
		logarithm_table[280] = 10'b00011_00100;
		logarithm_table[281] = 10'b00011_00100;
		logarithm_table[282] = 10'b00011_00100;
		logarithm_table[283] = 10'b00011_00101;
		logarithm_table[284] = 10'b00011_00101;
		logarithm_table[285] = 10'b00011_00101;
		logarithm_table[286] = 10'b00011_00101;
		logarithm_table[287] = 10'b00011_00101;
		logarithm_table[288] = 10'b00011_00101;
		logarithm_table[289] = 10'b00011_00110;
		logarithm_table[290] = 10'b00011_00110;
		logarithm_table[291] = 10'b00011_00110;
		logarithm_table[292] = 10'b00011_00110;
		logarithm_table[293] = 10'b00011_00110;
		logarithm_table[294] = 10'b00011_00110;
		logarithm_table[295] = 10'b00011_00111;
		logarithm_table[296] = 10'b00011_00111;
		logarithm_table[297] = 10'b00011_00111;
		logarithm_table[298] = 10'b00011_00111;
		logarithm_table[299] = 10'b00011_00111;
		logarithm_table[300] = 10'b00011_00111;
		logarithm_table[301] = 10'b00011_00111;
		logarithm_table[302] = 10'b00011_01000;
		logarithm_table[303] = 10'b00011_01000;
		logarithm_table[304] = 10'b00011_01000;
		logarithm_table[305] = 10'b00011_01000;
		logarithm_table[306] = 10'b00011_01000;
		logarithm_table[307] = 10'b00011_01000;
		logarithm_table[308] = 10'b00011_01001;
		logarithm_table[309] = 10'b00011_01001;
		logarithm_table[310] = 10'b00011_01001;
		logarithm_table[311] = 10'b00011_01001;
		logarithm_table[312] = 10'b00011_01001;
		logarithm_table[313] = 10'b00011_01001;
		logarithm_table[314] = 10'b00011_01001;
		logarithm_table[315] = 10'b00011_01010;
		logarithm_table[316] = 10'b00011_01010;
		logarithm_table[317] = 10'b00011_01010;
		logarithm_table[318] = 10'b00011_01010;
		logarithm_table[319] = 10'b00011_01010;
		logarithm_table[320] = 10'b00011_01010;
		logarithm_table[321] = 10'b00011_01010;
		logarithm_table[322] = 10'b00011_01011;
		logarithm_table[323] = 10'b00011_01011;
		logarithm_table[324] = 10'b00011_01011;
		logarithm_table[325] = 10'b00011_01011;
		logarithm_table[326] = 10'b00011_01011;
		logarithm_table[327] = 10'b00011_01011;
		logarithm_table[328] = 10'b00011_01011;
		logarithm_table[329] = 10'b00011_01100;
		logarithm_table[330] = 10'b00011_01100;
		logarithm_table[331] = 10'b00011_01100;
		logarithm_table[332] = 10'b00011_01100;
		logarithm_table[333] = 10'b00011_01100;
		logarithm_table[334] = 10'b00011_01100;
		logarithm_table[335] = 10'b00011_01100;
		logarithm_table[336] = 10'b00011_01101;
		logarithm_table[337] = 10'b00011_01101;
		logarithm_table[338] = 10'b00011_01101;
		logarithm_table[339] = 10'b00011_01101;
		logarithm_table[340] = 10'b00011_01101;
		logarithm_table[341] = 10'b00011_01101;
		logarithm_table[342] = 10'b00011_01101;
		logarithm_table[343] = 10'b00011_01110;
		logarithm_table[344] = 10'b00011_01110;
		logarithm_table[345] = 10'b00011_01110;
		logarithm_table[346] = 10'b00011_01110;
		logarithm_table[347] = 10'b00011_01110;
		logarithm_table[348] = 10'b00011_01110;
		logarithm_table[349] = 10'b00011_01110;
		logarithm_table[350] = 10'b00011_01110;
		logarithm_table[351] = 10'b00011_01111;
		logarithm_table[352] = 10'b00011_01111;
		logarithm_table[353] = 10'b00011_01111;
		logarithm_table[354] = 10'b00011_01111;
		logarithm_table[355] = 10'b00011_01111;
		logarithm_table[356] = 10'b00011_01111;
		logarithm_table[357] = 10'b00011_01111;
		logarithm_table[358] = 10'b00011_01111;
		logarithm_table[359] = 10'b00011_10000;
		logarithm_table[360] = 10'b00011_10000;
		logarithm_table[361] = 10'b00011_10000;
		logarithm_table[362] = 10'b00011_10000;
		logarithm_table[363] = 10'b00011_10000;
		logarithm_table[364] = 10'b00011_10000;
		logarithm_table[365] = 10'b00011_10000;
		logarithm_table[366] = 10'b00011_10001;
		logarithm_table[367] = 10'b00011_10001;
		logarithm_table[368] = 10'b00011_10001;
		logarithm_table[369] = 10'b00011_10001;
		logarithm_table[370] = 10'b00011_10001;
		logarithm_table[371] = 10'b00011_10001;
		logarithm_table[372] = 10'b00011_10001;
		logarithm_table[373] = 10'b00011_10001;
		logarithm_table[374] = 10'b00011_10010;
		logarithm_table[375] = 10'b00011_10010;
		logarithm_table[376] = 10'b00011_10010;
		logarithm_table[377] = 10'b00011_10010;
		logarithm_table[378] = 10'b00011_10010;
		logarithm_table[379] = 10'b00011_10010;
		logarithm_table[380] = 10'b00011_10010;
		logarithm_table[381] = 10'b00011_10010;
		logarithm_table[382] = 10'b00011_10010;
		logarithm_table[383] = 10'b00011_10011;
		logarithm_table[384] = 10'b00011_10011;
		logarithm_table[385] = 10'b00011_10011;
		logarithm_table[386] = 10'b00011_10011;
		logarithm_table[387] = 10'b00011_10011;
		logarithm_table[388] = 10'b00011_10011;
		logarithm_table[389] = 10'b00011_10011;
		logarithm_table[390] = 10'b00011_10011;
		logarithm_table[391] = 10'b00011_10100;
		logarithm_table[392] = 10'b00011_10100;
		logarithm_table[393] = 10'b00011_10100;
		logarithm_table[394] = 10'b00011_10100;
		logarithm_table[395] = 10'b00011_10100;
		logarithm_table[396] = 10'b00011_10100;
		logarithm_table[397] = 10'b00011_10100;
		logarithm_table[398] = 10'b00011_10100;
		logarithm_table[399] = 10'b00011_10100;
		logarithm_table[400] = 10'b00011_10101;
		logarithm_table[401] = 10'b00011_10101;
		logarithm_table[402] = 10'b00011_10101;
		logarithm_table[403] = 10'b00011_10101;
		logarithm_table[404] = 10'b00011_10101;
		logarithm_table[405] = 10'b00011_10101;
		logarithm_table[406] = 10'b00011_10101;
		logarithm_table[407] = 10'b00011_10101;
		logarithm_table[408] = 10'b00011_10110;
		logarithm_table[409] = 10'b00011_10110;
		logarithm_table[410] = 10'b00011_10110;
		logarithm_table[411] = 10'b00011_10110;
		logarithm_table[412] = 10'b00011_10110;
		logarithm_table[413] = 10'b00011_10110;
		logarithm_table[414] = 10'b00011_10110;
		logarithm_table[415] = 10'b00011_10110;
		logarithm_table[416] = 10'b00011_10110;
		logarithm_table[417] = 10'b00011_10111;
		logarithm_table[418] = 10'b00011_10111;
		logarithm_table[419] = 10'b00011_10111;
		logarithm_table[420] = 10'b00011_10111;
		logarithm_table[421] = 10'b00011_10111;
		logarithm_table[422] = 10'b00011_10111;
		logarithm_table[423] = 10'b00011_10111;
		logarithm_table[424] = 10'b00011_10111;
		logarithm_table[425] = 10'b00011_10111;
		logarithm_table[426] = 10'b00011_11000;
		logarithm_table[427] = 10'b00011_11000;
		logarithm_table[428] = 10'b00011_11000;
		logarithm_table[429] = 10'b00011_11000;
		logarithm_table[430] = 10'b00011_11000;
		logarithm_table[431] = 10'b00011_11000;
		logarithm_table[432] = 10'b00011_11000;
		logarithm_table[433] = 10'b00011_11000;
		logarithm_table[434] = 10'b00011_11000;
		logarithm_table[435] = 10'b00011_11000;
		logarithm_table[436] = 10'b00011_11001;
		logarithm_table[437] = 10'b00011_11001;
		logarithm_table[438] = 10'b00011_11001;
		logarithm_table[439] = 10'b00011_11001;
		logarithm_table[440] = 10'b00011_11001;
		logarithm_table[441] = 10'b00011_11001;
		logarithm_table[442] = 10'b00011_11001;
		logarithm_table[443] = 10'b00011_11001;
		logarithm_table[444] = 10'b00011_11001;
		logarithm_table[445] = 10'b00011_11010;
		logarithm_table[446] = 10'b00011_11010;
		logarithm_table[447] = 10'b00011_11010;
		logarithm_table[448] = 10'b00011_11010;
		logarithm_table[449] = 10'b00011_11010;
		logarithm_table[450] = 10'b00011_11010;
		logarithm_table[451] = 10'b00011_11010;
		logarithm_table[452] = 10'b00011_11010;
		logarithm_table[453] = 10'b00011_11010;
		logarithm_table[454] = 10'b00011_11010;
		logarithm_table[455] = 10'b00011_11011;
		logarithm_table[456] = 10'b00011_11011;
		logarithm_table[457] = 10'b00011_11011;
		logarithm_table[458] = 10'b00011_11011;
		logarithm_table[459] = 10'b00011_11011;
		logarithm_table[460] = 10'b00011_11011;
		logarithm_table[461] = 10'b00011_11011;
		logarithm_table[462] = 10'b00011_11011;
		logarithm_table[463] = 10'b00011_11011;
		logarithm_table[464] = 10'b00011_11011;
		logarithm_table[465] = 10'b00011_11100;
		logarithm_table[466] = 10'b00011_11100;
		logarithm_table[467] = 10'b00011_11100;
		logarithm_table[468] = 10'b00011_11100;
		logarithm_table[469] = 10'b00011_11100;
		logarithm_table[470] = 10'b00011_11100;
		logarithm_table[471] = 10'b00011_11100;
		logarithm_table[472] = 10'b00011_11100;
		logarithm_table[473] = 10'b00011_11100;
		logarithm_table[474] = 10'b00011_11100;
		logarithm_table[475] = 10'b00011_11101;
		logarithm_table[476] = 10'b00011_11101;
		logarithm_table[477] = 10'b00011_11101;
		logarithm_table[478] = 10'b00011_11101;
		logarithm_table[479] = 10'b00011_11101;
		logarithm_table[480] = 10'b00011_11101;
		logarithm_table[481] = 10'b00011_11101;
		logarithm_table[482] = 10'b00011_11101;
		logarithm_table[483] = 10'b00011_11101;
		logarithm_table[484] = 10'b00011_11101;
		logarithm_table[485] = 10'b00011_11101;
		logarithm_table[486] = 10'b00011_11110;
		logarithm_table[487] = 10'b00011_11110;
		logarithm_table[488] = 10'b00011_11110;
		logarithm_table[489] = 10'b00011_11110;
		logarithm_table[490] = 10'b00011_11110;
		logarithm_table[491] = 10'b00011_11110;
		logarithm_table[492] = 10'b00011_11110;
		logarithm_table[493] = 10'b00011_11110;
		logarithm_table[494] = 10'b00011_11110;
		logarithm_table[495] = 10'b00011_11110;
		logarithm_table[496] = 10'b00011_11111;
		logarithm_table[497] = 10'b00011_11111;
		logarithm_table[498] = 10'b00011_11111;
		logarithm_table[499] = 10'b00011_11111;
		logarithm_table[500] = 10'b00011_11111;
		logarithm_table[501] = 10'b00011_11111;
		logarithm_table[502] = 10'b00011_11111;
		logarithm_table[503] = 10'b00011_11111;
		logarithm_table[504] = 10'b00011_11111;
		logarithm_table[505] = 10'b00011_11111;
		logarithm_table[506] = 10'b00011_11111;
		logarithm_table[507] = 10'b00100_00000;
		logarithm_table[508] = 10'b00100_00000;
		logarithm_table[509] = 10'b00100_00000;
		logarithm_table[510] = 10'b00100_00000;
		logarithm_table[511] = 10'b00100_00000;
		Dminus[1] = 10'b11010_01111;
		Dminus[2] = 10'b11011_01110;
		Dminus[3] = 10'b11100_00000;
		Dminus[4] = 10'b11100_01101;
		Dminus[5] = 10'b11100_10111;
		Dminus[6] = 10'b11100_11111;
		Dminus[7] = 10'b11101_00101;
		Dminus[8] = 10'b11101_01011;
		Dminus[9] = 10'b11101_10000;
		Dminus[10] = 10'b11101_10100;
		Dminus[11] = 10'b11101_11000;
		Dminus[12] = 10'b11101_11100;
		Dminus[13] = 10'b11101_11111;
		Dminus[14] = 10'b11110_00010;
		Dminus[15] = 10'b11110_00101;
		Dminus[16] = 10'b11110_00111;
		Dminus[17] = 10'b11110_01010;
		Dminus[18] = 10'b11110_01100;
		Dminus[19] = 10'b11110_01110;
		Dminus[20] = 10'b11110_10000;
		Dminus[21] = 10'b11110_10010;
		Dminus[22] = 10'b11110_10011;
		Dminus[23] = 10'b11110_10101;
		Dminus[24] = 10'b11110_10110;
		Dminus[25] = 10'b11110_11000;
		Dminus[26] = 10'b11110_11001;
		Dminus[27] = 10'b11110_11010;
		Dminus[28] = 10'b11110_11100;
		Dminus[29] = 10'b11110_11101;
		Dminus[30] = 10'b11110_11110;
		Dminus[31] = 10'b11110_11111;
		Dminus[32] = 10'b11111_00000;
		Dminus[33] = 10'b11111_00001;
		Dminus[34] = 10'b11111_00010;
		Dminus[35] = 10'b11111_00011;
		Dminus[36] = 10'b11111_00100;
		Dminus[37] = 10'b11111_00101;
		Dminus[38] = 10'b11111_00101;
		Dminus[39] = 10'b11111_00110;
		Dminus[40] = 10'b11111_00111;
		Dminus[41] = 10'b11111_01000;
		Dminus[42] = 10'b11111_01000;
		Dminus[43] = 10'b11111_01001;
		Dminus[44] = 10'b11111_01010;
		Dminus[45] = 10'b11111_01010;
		Dminus[46] = 10'b11111_01011;
		Dminus[47] = 10'b11111_01011;
		Dminus[48] = 10'b11111_01100;
		Dminus[49] = 10'b11111_01100;
		Dminus[50] = 10'b11111_01101;
		Dminus[51] = 10'b11111_01101;
		Dminus[52] = 10'b11111_01110;
		Dminus[53] = 10'b11111_01110;
		Dminus[54] = 10'b11111_01111;
		Dminus[55] = 10'b11111_01111;
		Dminus[56] = 10'b11111_10000;
		Dminus[57] = 10'b11111_10000;
		Dminus[58] = 10'b11111_10001;
		Dminus[59] = 10'b11111_10001;
		Dminus[60] = 10'b11111_10001;
		Dminus[61] = 10'b11111_10010;
		Dminus[62] = 10'b11111_10010;
		Dminus[63] = 10'b11111_10010;
		Dminus[64] = 10'b11111_10011;
		Dminus[65] = 10'b11111_10011;
		Dminus[66] = 10'b11111_10011;
		Dminus[67] = 10'b11111_10100;
		Dminus[68] = 10'b11111_10100;
		Dminus[69] = 10'b11111_10100;
		Dminus[70] = 10'b11111_10101;
		Dminus[71] = 10'b11111_10101;
		Dminus[72] = 10'b11111_10101;
		Dminus[73] = 10'b11111_10101;
		Dminus[74] = 10'b11111_10110;
		Dminus[75] = 10'b11111_10110;
		Dminus[76] = 10'b11111_10110;
		Dminus[77] = 10'b11111_10110;
		Dminus[78] = 10'b11111_10111;
		Dminus[79] = 10'b11111_10111;
		Dminus[80] = 10'b11111_10111;
		Dminus[81] = 10'b11111_10111;
		Dminus[82] = 10'b11111_10111;
		Dminus[83] = 10'b11111_11000;
		Dminus[84] = 10'b11111_11000;
		Dminus[85] = 10'b11111_11000;
		Dminus[86] = 10'b11111_11000;
		Dminus[87] = 10'b11111_11000;
		Dminus[88] = 10'b11111_11001;
		Dminus[89] = 10'b11111_11001;
		Dminus[90] = 10'b11111_11001;
		Dminus[91] = 10'b11111_11001;
		Dminus[92] = 10'b11111_11001;
		Dminus[93] = 10'b11111_11001;
		Dminus[94] = 10'b11111_11010;
		Dminus[95] = 10'b11111_11010;
		Dminus[96] = 10'b11111_11010;
		Dminus[97] = 10'b11111_11010;
		Dminus[98] = 10'b11111_11010;
		Dminus[99] = 10'b11111_11010;
		Dminus[100] = 10'b11111_11010;
		Dminus[101] = 10'b11111_11011;
		Dminus[102] = 10'b11111_11011;
		Dminus[103] = 10'b11111_11011;
		Dminus[104] = 10'b11111_11011;
		Dminus[105] = 10'b11111_11011;
		Dminus[106] = 10'b11111_11011;
		Dminus[107] = 10'b11111_11011;
		Dminus[108] = 10'b11111_11011;
		Dminus[109] = 10'b11111_11011;
		Dminus[110] = 10'b11111_11100;
		Dminus[111] = 10'b11111_11100;
		Dminus[112] = 10'b11111_11100;
		Dminus[113] = 10'b11111_11100;
		Dminus[114] = 10'b11111_11100;
		Dminus[115] = 10'b11111_11100;
		Dminus[116] = 10'b11111_11100;
		Dminus[117] = 10'b11111_11100;
		Dminus[118] = 10'b11111_11100;
		Dminus[119] = 10'b11111_11100;
		Dminus[120] = 10'b11111_11100;
		Dminus[121] = 10'b11111_11101;
		Dminus[122] = 10'b11111_11101;
		Dminus[123] = 10'b11111_11101;
		Dminus[124] = 10'b11111_11101;
		Dminus[125] = 10'b11111_11101;
		Dminus[126] = 10'b11111_11101;
		Dminus[127] = 10'b11111_11101;
		Dminus[128] = 10'b11111_11101;
		Dminus[129] = 10'b11111_11101;
		Dminus[130] = 10'b11111_11101;
		Dminus[131] = 10'b11111_11101;
		Dminus[132] = 10'b11111_11101;
		Dminus[133] = 10'b11111_11101;
		Dminus[134] = 10'b11111_11101;
		Dminus[135] = 10'b11111_11101;
		Dminus[136] = 10'b11111_11110;
		Dminus[137] = 10'b11111_11110;
		Dminus[138] = 10'b11111_11110;
		Dminus[139] = 10'b11111_11110;
		Dminus[140] = 10'b11111_11110;
		Dminus[141] = 10'b11111_11110;
		Dminus[142] = 10'b11111_11110;
		Dminus[143] = 10'b11111_11110;
		Dminus[144] = 10'b11111_11110;
		Dminus[145] = 10'b11111_11110;
		Dminus[146] = 10'b11111_11110;
		Dminus[147] = 10'b11111_11110;
		Dminus[148] = 10'b11111_11110;
		Dminus[149] = 10'b11111_11110;
		Dminus[150] = 10'b11111_11110;
		Dminus[151] = 10'b11111_11110;
		Dminus[152] = 10'b11111_11110;
		Dminus[153] = 10'b11111_11110;
		Dminus[154] = 10'b11111_11110;
		Dminus[155] = 10'b11111_11110;
		Dminus[156] = 10'b11111_11110;
		Dminus[157] = 10'b11111_11110;
		Dminus[158] = 10'b11111_11110;
		Dminus[159] = 10'b11111_11111;
		Dminus[160] = 10'b11111_11111;
		Dminus[161] = 10'b11111_11111;
		Dminus[162] = 10'b11111_11111;
		Dminus[163] = 10'b11111_11111;
		Dminus[164] = 10'b11111_11111;
		Dminus[165] = 10'b11111_11111;
		Dminus[166] = 10'b11111_11111;
		Dminus[167] = 10'b11111_11111;
		Dminus[168] = 10'b11111_11111;
		Dminus[169] = 10'b11111_11111;
		Dminus[170] = 10'b11111_11111;
		Dminus[171] = 10'b11111_11111;
		Dminus[172] = 10'b11111_11111;
		Dminus[173] = 10'b11111_11111;
		Dminus[174] = 10'b11111_11111;
		Dminus[175] = 10'b11111_11111;
		Dminus[176] = 10'b11111_11111;
		Dminus[177] = 10'b11111_11111;
		Dminus[178] = 10'b11111_11111;
		Dminus[179] = 10'b11111_11111;
		Dminus[180] = 10'b11111_11111;
		Dminus[181] = 10'b11111_11111;
		Dminus[182] = 10'b11111_11111;
		Dminus[183] = 10'b11111_11111;
		Dminus[184] = 10'b11111_11111;
		Dminus[185] = 10'b11111_11111;
		Dminus[186] = 10'b11111_11111;
		Dminus[187] = 10'b11111_11111;
		Dminus[188] = 10'b11111_11111;
		Dminus[189] = 10'b11111_11111;
		Dminus[190] = 10'b11111_11111;
		Dminus[191] = 10'b11111_11111;
		Dminus[192] = 10'b11111_11111;
		Dminus[193] = 10'b11111_11111;
		Dminus[194] = 10'b11111_11111;
		Dminus[195] = 10'b11111_11111;
		Dminus[196] = 10'b11111_11111;
		Dminus[197] = 10'b11111_11111;
		Dminus[198] = 10'b11111_11111;
		Dminus[199] = 10'b11111_11111;
		Dminus[200] = 10'b11111_11111;
		Dminus[201] = 10'b11111_11111;
		Dminus[202] = 10'b11111_11111;
		Dminus[203] = 10'b11111_11111;
		Dminus[204] = 10'b11111_11111;
		Dminus[205] = 10'b11111_11111;
		Dminus[206] = 10'b11111_11111;
		Dminus[207] = 10'b11111_11111;
		Dminus[208] = 10'b11111_11111;
		Dminus[209] = 10'b11111_11111;
		Dminus[210] = 10'b00000_00000;
		Dminus[211] = 10'b00000_00000;
		Dminus[212] = 10'b00000_00000;
		Dminus[213] = 10'b00000_00000;
		Dminus[214] = 10'b00000_00000;
		Dminus[215] = 10'b00000_00000;
		Dminus[216] = 10'b00000_00000;
		Dminus[217] = 10'b00000_00000;
		Dminus[218] = 10'b00000_00000;
		Dminus[219] = 10'b00000_00000;
		Dminus[220] = 10'b00000_00000;
		Dminus[221] = 10'b00000_00000;
		Dminus[222] = 10'b00000_00000;
		Dminus[223] = 10'b00000_00000;
		Dminus[224] = 10'b00000_00000;
		Dminus[225] = 10'b00000_00000;
		Dminus[226] = 10'b00000_00000;
		Dminus[227] = 10'b00000_00000;
		Dminus[228] = 10'b00000_00000;
		Dminus[229] = 10'b00000_00000;
		Dminus[230] = 10'b00000_00000;
		Dminus[231] = 10'b00000_00000;
		Dminus[232] = 10'b00000_00000;
		Dminus[233] = 10'b00000_00000;
		Dminus[234] = 10'b00000_00000;
		Dminus[235] = 10'b00000_00000;
		Dminus[236] = 10'b00000_00000;
		Dminus[237] = 10'b00000_00000;
		Dminus[238] = 10'b00000_00000;
		Dminus[239] = 10'b00000_00000;
		Dminus[240] = 10'b00000_00000;
		Dminus[241] = 10'b00000_00000;
		Dminus[242] = 10'b00000_00000;
		Dminus[243] = 10'b00000_00000;
		Dminus[244] = 10'b00000_00000;
		Dminus[245] = 10'b00000_00000;
		Dminus[246] = 10'b00000_00000;
		Dminus[247] = 10'b00000_00000;
		Dminus[248] = 10'b00000_00000;
		Dminus[249] = 10'b00000_00000;
		Dminus[250] = 10'b00000_00000;
		Dminus[251] = 10'b00000_00000;
		Dminus[252] = 10'b00000_00000;
		Dminus[253] = 10'b00000_00000;
		Dminus[254] = 10'b00000_00000;
		Dminus[255] = 10'b00000_00000;
		Dminus[256] = 10'b00000_00000;
		Dminus[257] = 10'b00000_00000;
		Dminus[258] = 10'b00000_00000;
		Dminus[259] = 10'b00000_00000;
		Dminus[260] = 10'b00000_00000;
		Dminus[261] = 10'b00000_00000;
		Dminus[262] = 10'b00000_00000;
		Dminus[263] = 10'b00000_00000;
		Dminus[264] = 10'b00000_00000;
		Dminus[265] = 10'b00000_00000;
		Dminus[266] = 10'b00000_00000;
		Dminus[267] = 10'b00000_00000;
		Dminus[268] = 10'b00000_00000;
		Dminus[269] = 10'b00000_00000;
		Dminus[270] = 10'b00000_00000;
		Dminus[271] = 10'b00000_00000;
		Dminus[272] = 10'b00000_00000;
		Dminus[273] = 10'b00000_00000;
		Dminus[274] = 10'b00000_00000;
		Dminus[275] = 10'b00000_00000;
		Dminus[276] = 10'b00000_00000;
		Dminus[277] = 10'b00000_00000;
		Dminus[278] = 10'b00000_00000;
		Dminus[279] = 10'b00000_00000;
		Dminus[280] = 10'b00000_00000;
		Dminus[281] = 10'b00000_00000;
		Dminus[282] = 10'b00000_00000;
		Dminus[283] = 10'b00000_00000;
		Dminus[284] = 10'b00000_00000;
		Dminus[285] = 10'b00000_00000;
		Dminus[286] = 10'b00000_00000;
		Dminus[287] = 10'b00000_00000;
		Dminus[288] = 10'b00000_00000;
		Dminus[289] = 10'b00000_00000;
		Dminus[290] = 10'b00000_00000;
		Dminus[291] = 10'b00000_00000;
		Dminus[292] = 10'b00000_00000;
		Dminus[293] = 10'b00000_00000;
		Dminus[294] = 10'b00000_00000;
		Dminus[295] = 10'b00000_00000;
		Dminus[296] = 10'b00000_00000;
		Dminus[297] = 10'b00000_00000;
		Dminus[298] = 10'b00000_00000;
		Dminus[299] = 10'b00000_00000;
		Dminus[300] = 10'b00000_00000;
		Dminus[301] = 10'b00000_00000;
		Dminus[302] = 10'b00000_00000;
		Dminus[303] = 10'b00000_00000;
		Dminus[304] = 10'b00000_00000;
		Dminus[305] = 10'b00000_00000;
		Dminus[306] = 10'b00000_00000;
		Dminus[307] = 10'b00000_00000;
		Dminus[308] = 10'b00000_00000;
		Dminus[309] = 10'b00000_00000;
		Dminus[310] = 10'b00000_00000;
		Dminus[311] = 10'b00000_00000;
		Dminus[312] = 10'b00000_00000;
		Dminus[313] = 10'b00000_00000;
		Dminus[314] = 10'b00000_00000;
		Dminus[315] = 10'b00000_00000;
		Dminus[316] = 10'b00000_00000;
		Dminus[317] = 10'b00000_00000;
		Dminus[318] = 10'b00000_00000;
		Dminus[319] = 10'b00000_00000;
		Dminus[320] = 10'b00000_00000;
		Dminus[321] = 10'b00000_00000;
		Dminus[322] = 10'b00000_00000;
		Dminus[323] = 10'b00000_00000;
		Dminus[324] = 10'b00000_00000;
		Dminus[325] = 10'b00000_00000;
		Dminus[326] = 10'b00000_00000;
		Dminus[327] = 10'b00000_00000;
		Dminus[328] = 10'b00000_00000;
		Dminus[329] = 10'b00000_00000;
		Dminus[330] = 10'b00000_00000;
		Dminus[331] = 10'b00000_00000;
		Dminus[332] = 10'b00000_00000;
		Dminus[333] = 10'b00000_00000;
		Dminus[334] = 10'b00000_00000;
		Dminus[335] = 10'b00000_00000;
		Dminus[336] = 10'b00000_00000;
		Dminus[337] = 10'b00000_00000;
		Dminus[338] = 10'b00000_00000;
		Dminus[339] = 10'b00000_00000;
		Dminus[340] = 10'b00000_00000;
		Dminus[341] = 10'b00000_00000;
		Dminus[342] = 10'b00000_00000;
		Dminus[343] = 10'b00000_00000;
		Dminus[344] = 10'b00000_00000;
		Dminus[345] = 10'b00000_00000;
		Dminus[346] = 10'b00000_00000;
		Dminus[347] = 10'b00000_00000;
		Dminus[348] = 10'b00000_00000;
		Dminus[349] = 10'b00000_00000;
		Dminus[350] = 10'b00000_00000;
		Dminus[351] = 10'b00000_00000;
		Dminus[352] = 10'b00000_00000;
		Dminus[353] = 10'b00000_00000;
		Dminus[354] = 10'b00000_00000;
		Dminus[355] = 10'b00000_00000;
		Dminus[356] = 10'b00000_00000;
		Dminus[357] = 10'b00000_00000;
		Dminus[358] = 10'b00000_00000;
		Dminus[359] = 10'b00000_00000;
		Dminus[360] = 10'b00000_00000;
		Dminus[361] = 10'b00000_00000;
		Dminus[362] = 10'b00000_00000;
		Dminus[363] = 10'b00000_00000;
		Dminus[364] = 10'b00000_00000;
		Dminus[365] = 10'b00000_00000;
		Dminus[366] = 10'b00000_00000;
		Dminus[367] = 10'b00000_00000;
		Dminus[368] = 10'b00000_00000;
		Dminus[369] = 10'b00000_00000;
		Dminus[370] = 10'b00000_00000;
		Dminus[371] = 10'b00000_00000;
		Dminus[372] = 10'b00000_00000;
		Dminus[373] = 10'b00000_00000;
		Dminus[374] = 10'b00000_00000;
		Dminus[375] = 10'b00000_00000;
		Dminus[376] = 10'b00000_00000;
		Dminus[377] = 10'b00000_00000;
		Dminus[378] = 10'b00000_00000;
		Dminus[379] = 10'b00000_00000;
		Dminus[380] = 10'b00000_00000;
		Dminus[381] = 10'b00000_00000;
		Dminus[382] = 10'b00000_00000;
		Dminus[383] = 10'b00000_00000;
		Dminus[384] = 10'b00000_00000;
		Dminus[385] = 10'b00000_00000;
		Dminus[386] = 10'b00000_00000;
		Dminus[387] = 10'b00000_00000;
		Dminus[388] = 10'b00000_00000;
		Dminus[389] = 10'b00000_00000;
		Dminus[390] = 10'b00000_00000;
		Dminus[391] = 10'b00000_00000;
		Dminus[392] = 10'b00000_00000;
		Dminus[393] = 10'b00000_00000;
		Dminus[394] = 10'b00000_00000;
		Dminus[395] = 10'b00000_00000;
		Dminus[396] = 10'b00000_00000;
		Dminus[397] = 10'b00000_00000;
		Dminus[398] = 10'b00000_00000;
		Dminus[399] = 10'b00000_00000;
		Dminus[400] = 10'b00000_00000;
		Dminus[401] = 10'b00000_00000;
		Dminus[402] = 10'b00000_00000;
		Dminus[403] = 10'b00000_00000;
		Dminus[404] = 10'b00000_00000;
		Dminus[405] = 10'b00000_00000;
		Dminus[406] = 10'b00000_00000;
		Dminus[407] = 10'b00000_00000;
		Dminus[408] = 10'b00000_00000;
		Dminus[409] = 10'b00000_00000;
		Dminus[410] = 10'b00000_00000;
		Dminus[411] = 10'b00000_00000;
		Dminus[412] = 10'b00000_00000;
		Dminus[413] = 10'b00000_00000;
		Dminus[414] = 10'b00000_00000;
		Dminus[415] = 10'b00000_00000;
		Dminus[416] = 10'b00000_00000;
		Dminus[417] = 10'b00000_00000;
		Dminus[418] = 10'b00000_00000;
		Dminus[419] = 10'b00000_00000;
		Dminus[420] = 10'b00000_00000;
		Dminus[421] = 10'b00000_00000;
		Dminus[422] = 10'b00000_00000;
		Dminus[423] = 10'b00000_00000;
		Dminus[424] = 10'b00000_00000;
		Dminus[425] = 10'b00000_00000;
		Dminus[426] = 10'b00000_00000;
		Dminus[427] = 10'b00000_00000;
		Dminus[428] = 10'b00000_00000;
		Dminus[429] = 10'b00000_00000;
		Dminus[430] = 10'b00000_00000;
		Dminus[431] = 10'b00000_00000;
		Dminus[432] = 10'b00000_00000;
		Dminus[433] = 10'b00000_00000;
		Dminus[434] = 10'b00000_00000;
		Dminus[435] = 10'b00000_00000;
		Dminus[436] = 10'b00000_00000;
		Dminus[437] = 10'b00000_00000;
		Dminus[438] = 10'b00000_00000;
		Dminus[439] = 10'b00000_00000;
		Dminus[440] = 10'b00000_00000;
		Dminus[441] = 10'b00000_00000;
		Dminus[442] = 10'b00000_00000;
		Dminus[443] = 10'b00000_00000;
		Dminus[444] = 10'b00000_00000;
		Dminus[445] = 10'b00000_00000;
		Dminus[446] = 10'b00000_00000;
		Dminus[447] = 10'b00000_00000;
		Dminus[448] = 10'b00000_00000;
		Dminus[449] = 10'b00000_00000;
		Dminus[450] = 10'b00000_00000;
		Dminus[451] = 10'b00000_00000;
		Dminus[452] = 10'b00000_00000;
		Dminus[453] = 10'b00000_00000;
		Dminus[454] = 10'b00000_00000;
		Dminus[455] = 10'b00000_00000;
		Dminus[456] = 10'b00000_00000;
		Dminus[457] = 10'b00000_00000;
		Dminus[458] = 10'b00000_00000;
		Dminus[459] = 10'b00000_00000;
		Dminus[460] = 10'b00000_00000;
		Dminus[461] = 10'b00000_00000;
		Dminus[462] = 10'b00000_00000;
		Dminus[463] = 10'b00000_00000;
		Dminus[464] = 10'b00000_00000;
		Dminus[465] = 10'b00000_00000;
		Dminus[466] = 10'b00000_00000;
		Dminus[467] = 10'b00000_00000;
		Dminus[468] = 10'b00000_00000;
		Dminus[469] = 10'b00000_00000;
		Dminus[470] = 10'b00000_00000;
		Dminus[471] = 10'b00000_00000;
		Dminus[472] = 10'b00000_00000;
		Dminus[473] = 10'b00000_00000;
		Dminus[474] = 10'b00000_00000;
		Dminus[475] = 10'b00000_00000;
		Dminus[476] = 10'b00000_00000;
		Dminus[477] = 10'b00000_00000;
		Dminus[478] = 10'b00000_00000;
		Dminus[479] = 10'b00000_00000;
		Dminus[480] = 10'b00000_00000;
		Dminus[481] = 10'b00000_00000;
		Dminus[482] = 10'b00000_00000;
		Dminus[483] = 10'b00000_00000;
		Dminus[484] = 10'b00000_00000;
		Dminus[485] = 10'b00000_00000;
		Dminus[486] = 10'b00000_00000;
		Dminus[487] = 10'b00000_00000;
		Dminus[488] = 10'b00000_00000;
		Dminus[489] = 10'b00000_00000;
		Dminus[490] = 10'b00000_00000;
		Dminus[491] = 10'b00000_00000;
		Dminus[492] = 10'b00000_00000;
		Dminus[493] = 10'b00000_00000;
		Dminus[494] = 10'b00000_00000;
		Dminus[495] = 10'b00000_00000;
		Dminus[496] = 10'b00000_00000;
		Dminus[497] = 10'b00000_00000;
		Dminus[498] = 10'b00000_00000;
		Dminus[499] = 10'b00000_00000;
		Dminus[500] = 10'b00000_00000;
		Dminus[501] = 10'b00000_00000;
		Dminus[502] = 10'b00000_00000;
		Dminus[503] = 10'b00000_00000;
		Dminus[504] = 10'b00000_00000;
		Dminus[505] = 10'b00000_00000;
		Dminus[506] = 10'b00000_00000;
		Dminus[507] = 10'b00000_00000;
		Dminus[508] = 10'b00000_00000;
		Dminus[509] = 10'b00000_00000;
		Dminus[510] = 10'b00000_00000;
		Dminus[511] = 10'b00000_00000;
		Dplus[1] = 10'b00001_00000;
		Dplus[2] = 10'b00000_11111;
		Dplus[3] = 10'b00000_11111;
		Dplus[4] = 10'b00000_11110;
		Dplus[5] = 10'b00000_11110;
		Dplus[6] = 10'b00000_11101;
		Dplus[7] = 10'b00000_11101;
		Dplus[8] = 10'b00000_11100;
		Dplus[9] = 10'b00000_11100;
		Dplus[10] = 10'b00000_11011;
		Dplus[11] = 10'b00000_11011;
		Dplus[12] = 10'b00000_11010;
		Dplus[13] = 10'b00000_11010;
		Dplus[14] = 10'b00000_11010;
		Dplus[15] = 10'b00000_11001;
		Dplus[16] = 10'b00000_11001;
		Dplus[17] = 10'b00000_11000;
		Dplus[18] = 10'b00000_11000;
		Dplus[19] = 10'b00000_10111;
		Dplus[20] = 10'b00000_10111;
		Dplus[21] = 10'b00000_10111;
		Dplus[22] = 10'b00000_10110;
		Dplus[23] = 10'b00000_10110;
		Dplus[24] = 10'b00000_10110;
		Dplus[25] = 10'b00000_10101;
		Dplus[26] = 10'b00000_10101;
		Dplus[27] = 10'b00000_10100;
		Dplus[28] = 10'b00000_10100;
		Dplus[29] = 10'b00000_10100;
		Dplus[30] = 10'b00000_10011;
		Dplus[31] = 10'b00000_10011;
		Dplus[32] = 10'b00000_10011;
		Dplus[33] = 10'b00000_10010;
		Dplus[34] = 10'b00000_10010;
		Dplus[35] = 10'b00000_10010;
		Dplus[36] = 10'b00000_10001;
		Dplus[37] = 10'b00000_10001;
		Dplus[38] = 10'b00000_10001;
		Dplus[39] = 10'b00000_10001;
		Dplus[40] = 10'b00000_10000;
		Dplus[41] = 10'b00000_10000;
		Dplus[42] = 10'b00000_10000;
		Dplus[43] = 10'b00000_01111;
		Dplus[44] = 10'b00000_01111;
		Dplus[45] = 10'b00000_01111;
		Dplus[46] = 10'b00000_01111;
		Dplus[47] = 10'b00000_01110;
		Dplus[48] = 10'b00000_01110;
		Dplus[49] = 10'b00000_01110;
		Dplus[50] = 10'b00000_01101;
		Dplus[51] = 10'b00000_01101;
		Dplus[52] = 10'b00000_01101;
		Dplus[53] = 10'b00000_01101;
		Dplus[54] = 10'b00000_01100;
		Dplus[55] = 10'b00000_01100;
		Dplus[56] = 10'b00000_01100;
		Dplus[57] = 10'b00000_01100;
		Dplus[58] = 10'b00000_01100;
		Dplus[59] = 10'b00000_01011;
		Dplus[60] = 10'b00000_01011;
		Dplus[61] = 10'b00000_01011;
		Dplus[62] = 10'b00000_01011;
		Dplus[63] = 10'b00000_01011;
		Dplus[64] = 10'b00000_01010;
		Dplus[65] = 10'b00000_01010;
		Dplus[66] = 10'b00000_01010;
		Dplus[67] = 10'b00000_01010;
		Dplus[68] = 10'b00000_01010;
		Dplus[69] = 10'b00000_01001;
		Dplus[70] = 10'b00000_01001;
		Dplus[71] = 10'b00000_01001;
		Dplus[72] = 10'b00000_01001;
		Dplus[73] = 10'b00000_01001;
		Dplus[74] = 10'b00000_01000;
		Dplus[75] = 10'b00000_01000;
		Dplus[76] = 10'b00000_01000;
		Dplus[77] = 10'b00000_01000;
		Dplus[78] = 10'b00000_01000;
		Dplus[79] = 10'b00000_01000;
		Dplus[80] = 10'b00000_01000;
		Dplus[81] = 10'b00000_00111;
		Dplus[82] = 10'b00000_00111;
		Dplus[83] = 10'b00000_00111;
		Dplus[84] = 10'b00000_00111;
		Dplus[85] = 10'b00000_00111;
		Dplus[86] = 10'b00000_00111;
		Dplus[87] = 10'b00000_00111;
		Dplus[88] = 10'b00000_00110;
		Dplus[89] = 10'b00000_00110;
		Dplus[90] = 10'b00000_00110;
		Dplus[91] = 10'b00000_00110;
		Dplus[92] = 10'b00000_00110;
		Dplus[93] = 10'b00000_00110;
		Dplus[94] = 10'b00000_00110;
		Dplus[95] = 10'b00000_00110;
		Dplus[96] = 10'b00000_00101;
		Dplus[97] = 10'b00000_00101;
		Dplus[98] = 10'b00000_00101;
		Dplus[99] = 10'b00000_00101;
		Dplus[100] = 10'b00000_00101;
		Dplus[101] = 10'b00000_00101;
		Dplus[102] = 10'b00000_00101;
		Dplus[103] = 10'b00000_00101;
		Dplus[104] = 10'b00000_00101;
		Dplus[105] = 10'b00000_00101;
		Dplus[106] = 10'b00000_00100;
		Dplus[107] = 10'b00000_00100;
		Dplus[108] = 10'b00000_00100;
		Dplus[109] = 10'b00000_00100;
		Dplus[110] = 10'b00000_00100;
		Dplus[111] = 10'b00000_00100;
		Dplus[112] = 10'b00000_00100;
		Dplus[113] = 10'b00000_00100;
		Dplus[114] = 10'b00000_00100;
		Dplus[115] = 10'b00000_00100;
		Dplus[116] = 10'b00000_00100;
		Dplus[117] = 10'b00000_00100;
		Dplus[118] = 10'b00000_00011;
		Dplus[119] = 10'b00000_00011;
		Dplus[120] = 10'b00000_00011;
		Dplus[121] = 10'b00000_00011;
		Dplus[122] = 10'b00000_00011;
		Dplus[123] = 10'b00000_00011;
		Dplus[124] = 10'b00000_00011;
		Dplus[125] = 10'b00000_00011;
		Dplus[126] = 10'b00000_00011;
		Dplus[127] = 10'b00000_00011;
		Dplus[128] = 10'b00000_00011;
		Dplus[129] = 10'b00000_00011;
		Dplus[130] = 10'b00000_00011;
		Dplus[131] = 10'b00000_00011;
		Dplus[132] = 10'b00000_00011;
		Dplus[133] = 10'b00000_00011;
		Dplus[134] = 10'b00000_00010;
		Dplus[135] = 10'b00000_00010;
		Dplus[136] = 10'b00000_00010;
		Dplus[137] = 10'b00000_00010;
		Dplus[138] = 10'b00000_00010;
		Dplus[139] = 10'b00000_00010;
		Dplus[140] = 10'b00000_00010;
		Dplus[141] = 10'b00000_00010;
		Dplus[142] = 10'b00000_00010;
		Dplus[143] = 10'b00000_00010;
		Dplus[144] = 10'b00000_00010;
		Dplus[145] = 10'b00000_00010;
		Dplus[146] = 10'b00000_00010;
		Dplus[147] = 10'b00000_00010;
		Dplus[148] = 10'b00000_00010;
		Dplus[149] = 10'b00000_00010;
		Dplus[150] = 10'b00000_00010;
		Dplus[151] = 10'b00000_00010;
		Dplus[152] = 10'b00000_00010;
		Dplus[153] = 10'b00000_00010;
		Dplus[154] = 10'b00000_00010;
		Dplus[155] = 10'b00000_00010;
		Dplus[156] = 10'b00000_00010;
		Dplus[157] = 10'b00000_00010;
		Dplus[158] = 10'b00000_00001;
		Dplus[159] = 10'b00000_00001;
		Dplus[160] = 10'b00000_00001;
		Dplus[161] = 10'b00000_00001;
		Dplus[162] = 10'b00000_00001;
		Dplus[163] = 10'b00000_00001;
		Dplus[164] = 10'b00000_00001;
		Dplus[165] = 10'b00000_00001;
		Dplus[166] = 10'b00000_00001;
		Dplus[167] = 10'b00000_00001;
		Dplus[168] = 10'b00000_00001;
		Dplus[169] = 10'b00000_00001;
		Dplus[170] = 10'b00000_00001;
		Dplus[171] = 10'b00000_00001;
		Dplus[172] = 10'b00000_00001;
		Dplus[173] = 10'b00000_00001;
		Dplus[174] = 10'b00000_00001;
		Dplus[175] = 10'b00000_00001;
		Dplus[176] = 10'b00000_00001;
		Dplus[177] = 10'b00000_00001;
		Dplus[178] = 10'b00000_00001;
		Dplus[179] = 10'b00000_00001;
		Dplus[180] = 10'b00000_00001;
		Dplus[181] = 10'b00000_00001;
		Dplus[182] = 10'b00000_00001;
		Dplus[183] = 10'b00000_00001;
		Dplus[184] = 10'b00000_00001;
		Dplus[185] = 10'b00000_00001;
		Dplus[186] = 10'b00000_00001;
		Dplus[187] = 10'b00000_00001;
		Dplus[188] = 10'b00000_00001;
		Dplus[189] = 10'b00000_00001;
		Dplus[190] = 10'b00000_00001;
		Dplus[191] = 10'b00000_00001;
		Dplus[192] = 10'b00000_00001;
		Dplus[193] = 10'b00000_00001;
		Dplus[194] = 10'b00000_00001;
		Dplus[195] = 10'b00000_00001;
		Dplus[196] = 10'b00000_00001;
		Dplus[197] = 10'b00000_00001;
		Dplus[198] = 10'b00000_00001;
		Dplus[199] = 10'b00000_00001;
		Dplus[200] = 10'b00000_00001;
		Dplus[201] = 10'b00000_00001;
		Dplus[202] = 10'b00000_00001;
		Dplus[203] = 10'b00000_00001;
		Dplus[204] = 10'b00000_00001;
		Dplus[205] = 10'b00000_00001;
		Dplus[206] = 10'b00000_00001;
		Dplus[207] = 10'b00000_00001;
		Dplus[208] = 10'b00000_00001;
		Dplus[209] = 10'b00000_00000;
		Dplus[210] = 10'b00000_00000;
		Dplus[211] = 10'b00000_00000;
		Dplus[212] = 10'b00000_00000;
		Dplus[213] = 10'b00000_00000;
		Dplus[214] = 10'b00000_00000;
		Dplus[215] = 10'b00000_00000;
		Dplus[216] = 10'b00000_00000;
		Dplus[217] = 10'b00000_00000;
		Dplus[218] = 10'b00000_00000;
		Dplus[219] = 10'b00000_00000;
		Dplus[220] = 10'b00000_00000;
		Dplus[221] = 10'b00000_00000;
		Dplus[222] = 10'b00000_00000;
		Dplus[223] = 10'b00000_00000;
		Dplus[224] = 10'b00000_00000;
		Dplus[225] = 10'b00000_00000;
		Dplus[226] = 10'b00000_00000;
		Dplus[227] = 10'b00000_00000;
		Dplus[228] = 10'b00000_00000;
		Dplus[229] = 10'b00000_00000;
		Dplus[230] = 10'b00000_00000;
		Dplus[231] = 10'b00000_00000;
		Dplus[232] = 10'b00000_00000;
		Dplus[233] = 10'b00000_00000;
		Dplus[234] = 10'b00000_00000;
		Dplus[235] = 10'b00000_00000;
		Dplus[236] = 10'b00000_00000;
		Dplus[237] = 10'b00000_00000;
		Dplus[238] = 10'b00000_00000;
		Dplus[239] = 10'b00000_00000;
		Dplus[240] = 10'b00000_00000;
		Dplus[241] = 10'b00000_00000;
		Dplus[242] = 10'b00000_00000;
		Dplus[243] = 10'b00000_00000;
		Dplus[244] = 10'b00000_00000;
		Dplus[245] = 10'b00000_00000;
		Dplus[246] = 10'b00000_00000;
		Dplus[247] = 10'b00000_00000;
		Dplus[248] = 10'b00000_00000;
		Dplus[249] = 10'b00000_00000;
		Dplus[250] = 10'b00000_00000;
		Dplus[251] = 10'b00000_00000;
		Dplus[252] = 10'b00000_00000;
		Dplus[253] = 10'b00000_00000;
		Dplus[254] = 10'b00000_00000;
		Dplus[255] = 10'b00000_00000;
		Dplus[256] = 10'b00000_00000;
		Dplus[257] = 10'b00000_00000;
		Dplus[258] = 10'b00000_00000;
		Dplus[259] = 10'b00000_00000;
		Dplus[260] = 10'b00000_00000;
		Dplus[261] = 10'b00000_00000;
		Dplus[262] = 10'b00000_00000;
		Dplus[263] = 10'b00000_00000;
		Dplus[264] = 10'b00000_00000;
		Dplus[265] = 10'b00000_00000;
		Dplus[266] = 10'b00000_00000;
		Dplus[267] = 10'b00000_00000;
		Dplus[268] = 10'b00000_00000;
		Dplus[269] = 10'b00000_00000;
		Dplus[270] = 10'b00000_00000;
		Dplus[271] = 10'b00000_00000;
		Dplus[272] = 10'b00000_00000;
		Dplus[273] = 10'b00000_00000;
		Dplus[274] = 10'b00000_00000;
		Dplus[275] = 10'b00000_00000;
		Dplus[276] = 10'b00000_00000;
		Dplus[277] = 10'b00000_00000;
		Dplus[278] = 10'b00000_00000;
		Dplus[279] = 10'b00000_00000;
		Dplus[280] = 10'b00000_00000;
		Dplus[281] = 10'b00000_00000;
		Dplus[282] = 10'b00000_00000;
		Dplus[283] = 10'b00000_00000;
		Dplus[284] = 10'b00000_00000;
		Dplus[285] = 10'b00000_00000;
		Dplus[286] = 10'b00000_00000;
		Dplus[287] = 10'b00000_00000;
		Dplus[288] = 10'b00000_00000;
		Dplus[289] = 10'b00000_00000;
		Dplus[290] = 10'b00000_00000;
		Dplus[291] = 10'b00000_00000;
		Dplus[292] = 10'b00000_00000;
		Dplus[293] = 10'b00000_00000;
		Dplus[294] = 10'b00000_00000;
		Dplus[295] = 10'b00000_00000;
		Dplus[296] = 10'b00000_00000;
		Dplus[297] = 10'b00000_00000;
		Dplus[298] = 10'b00000_00000;
		Dplus[299] = 10'b00000_00000;
		Dplus[300] = 10'b00000_00000;
		Dplus[301] = 10'b00000_00000;
		Dplus[302] = 10'b00000_00000;
		Dplus[303] = 10'b00000_00000;
		Dplus[304] = 10'b00000_00000;
		Dplus[305] = 10'b00000_00000;
		Dplus[306] = 10'b00000_00000;
		Dplus[307] = 10'b00000_00000;
		Dplus[308] = 10'b00000_00000;
		Dplus[309] = 10'b00000_00000;
		Dplus[310] = 10'b00000_00000;
		Dplus[311] = 10'b00000_00000;
		Dplus[312] = 10'b00000_00000;
		Dplus[313] = 10'b00000_00000;
		Dplus[314] = 10'b00000_00000;
		Dplus[315] = 10'b00000_00000;
		Dplus[316] = 10'b00000_00000;
		Dplus[317] = 10'b00000_00000;
		Dplus[318] = 10'b00000_00000;
		Dplus[319] = 10'b00000_00000;
		Dplus[320] = 10'b00000_00000;
		Dplus[321] = 10'b00000_00000;
		Dplus[322] = 10'b00000_00000;
		Dplus[323] = 10'b00000_00000;
		Dplus[324] = 10'b00000_00000;
		Dplus[325] = 10'b00000_00000;
		Dplus[326] = 10'b00000_00000;
		Dplus[327] = 10'b00000_00000;
		Dplus[328] = 10'b00000_00000;
		Dplus[329] = 10'b00000_00000;
		Dplus[330] = 10'b00000_00000;
		Dplus[331] = 10'b00000_00000;
		Dplus[332] = 10'b00000_00000;
		Dplus[333] = 10'b00000_00000;
		Dplus[334] = 10'b00000_00000;
		Dplus[335] = 10'b00000_00000;
		Dplus[336] = 10'b00000_00000;
		Dplus[337] = 10'b00000_00000;
		Dplus[338] = 10'b00000_00000;
		Dplus[339] = 10'b00000_00000;
		Dplus[340] = 10'b00000_00000;
		Dplus[341] = 10'b00000_00000;
		Dplus[342] = 10'b00000_00000;
		Dplus[343] = 10'b00000_00000;
		Dplus[344] = 10'b00000_00000;
		Dplus[345] = 10'b00000_00000;
		Dplus[346] = 10'b00000_00000;
		Dplus[347] = 10'b00000_00000;
		Dplus[348] = 10'b00000_00000;
		Dplus[349] = 10'b00000_00000;
		Dplus[350] = 10'b00000_00000;
		Dplus[351] = 10'b00000_00000;
		Dplus[352] = 10'b00000_00000;
		Dplus[353] = 10'b00000_00000;
		Dplus[354] = 10'b00000_00000;
		Dplus[355] = 10'b00000_00000;
		Dplus[356] = 10'b00000_00000;
		Dplus[357] = 10'b00000_00000;
		Dplus[358] = 10'b00000_00000;
		Dplus[359] = 10'b00000_00000;
		Dplus[360] = 10'b00000_00000;
		Dplus[361] = 10'b00000_00000;
		Dplus[362] = 10'b00000_00000;
		Dplus[363] = 10'b00000_00000;
		Dplus[364] = 10'b00000_00000;
		Dplus[365] = 10'b00000_00000;
		Dplus[366] = 10'b00000_00000;
		Dplus[367] = 10'b00000_00000;
		Dplus[368] = 10'b00000_00000;
		Dplus[369] = 10'b00000_00000;
		Dplus[370] = 10'b00000_00000;
		Dplus[371] = 10'b00000_00000;
		Dplus[372] = 10'b00000_00000;
		Dplus[373] = 10'b00000_00000;
		Dplus[374] = 10'b00000_00000;
		Dplus[375] = 10'b00000_00000;
		Dplus[376] = 10'b00000_00000;
		Dplus[377] = 10'b00000_00000;
		Dplus[378] = 10'b00000_00000;
		Dplus[379] = 10'b00000_00000;
		Dplus[380] = 10'b00000_00000;
		Dplus[381] = 10'b00000_00000;
		Dplus[382] = 10'b00000_00000;
		Dplus[383] = 10'b00000_00000;
		Dplus[384] = 10'b00000_00000;
		Dplus[385] = 10'b00000_00000;
		Dplus[386] = 10'b00000_00000;
		Dplus[387] = 10'b00000_00000;
		Dplus[388] = 10'b00000_00000;
		Dplus[389] = 10'b00000_00000;
		Dplus[390] = 10'b00000_00000;
		Dplus[391] = 10'b00000_00000;
		Dplus[392] = 10'b00000_00000;
		Dplus[393] = 10'b00000_00000;
		Dplus[394] = 10'b00000_00000;
		Dplus[395] = 10'b00000_00000;
		Dplus[396] = 10'b00000_00000;
		Dplus[397] = 10'b00000_00000;
		Dplus[398] = 10'b00000_00000;
		Dplus[399] = 10'b00000_00000;
		Dplus[400] = 10'b00000_00000;
		Dplus[401] = 10'b00000_00000;
		Dplus[402] = 10'b00000_00000;
		Dplus[403] = 10'b00000_00000;
		Dplus[404] = 10'b00000_00000;
		Dplus[405] = 10'b00000_00000;
		Dplus[406] = 10'b00000_00000;
		Dplus[407] = 10'b00000_00000;
		Dplus[408] = 10'b00000_00000;
		Dplus[409] = 10'b00000_00000;
		Dplus[410] = 10'b00000_00000;
		Dplus[411] = 10'b00000_00000;
		Dplus[412] = 10'b00000_00000;
		Dplus[413] = 10'b00000_00000;
		Dplus[414] = 10'b00000_00000;
		Dplus[415] = 10'b00000_00000;
		Dplus[416] = 10'b00000_00000;
		Dplus[417] = 10'b00000_00000;
		Dplus[418] = 10'b00000_00000;
		Dplus[419] = 10'b00000_00000;
		Dplus[420] = 10'b00000_00000;
		Dplus[421] = 10'b00000_00000;
		Dplus[422] = 10'b00000_00000;
		Dplus[423] = 10'b00000_00000;
		Dplus[424] = 10'b00000_00000;
		Dplus[425] = 10'b00000_00000;
		Dplus[426] = 10'b00000_00000;
		Dplus[427] = 10'b00000_00000;
		Dplus[428] = 10'b00000_00000;
		Dplus[429] = 10'b00000_00000;
		Dplus[430] = 10'b00000_00000;
		Dplus[431] = 10'b00000_00000;
		Dplus[432] = 10'b00000_00000;
		Dplus[433] = 10'b00000_00000;
		Dplus[434] = 10'b00000_00000;
		Dplus[435] = 10'b00000_00000;
		Dplus[436] = 10'b00000_00000;
		Dplus[437] = 10'b00000_00000;
		Dplus[438] = 10'b00000_00000;
		Dplus[439] = 10'b00000_00000;
		Dplus[440] = 10'b00000_00000;
		Dplus[441] = 10'b00000_00000;
		Dplus[442] = 10'b00000_00000;
		Dplus[443] = 10'b00000_00000;
		Dplus[444] = 10'b00000_00000;
		Dplus[445] = 10'b00000_00000;
		Dplus[446] = 10'b00000_00000;
		Dplus[447] = 10'b00000_00000;
		Dplus[448] = 10'b00000_00000;
		Dplus[449] = 10'b00000_00000;
		Dplus[450] = 10'b00000_00000;
		Dplus[451] = 10'b00000_00000;
		Dplus[452] = 10'b00000_00000;
		Dplus[453] = 10'b00000_00000;
		Dplus[454] = 10'b00000_00000;
		Dplus[455] = 10'b00000_00000;
		Dplus[456] = 10'b00000_00000;
		Dplus[457] = 10'b00000_00000;
		Dplus[458] = 10'b00000_00000;
		Dplus[459] = 10'b00000_00000;
		Dplus[460] = 10'b00000_00000;
		Dplus[461] = 10'b00000_00000;
		Dplus[462] = 10'b00000_00000;
		Dplus[463] = 10'b00000_00000;
		Dplus[464] = 10'b00000_00000;
		Dplus[465] = 10'b00000_00000;
		Dplus[466] = 10'b00000_00000;
		Dplus[467] = 10'b00000_00000;
		Dplus[468] = 10'b00000_00000;
		Dplus[469] = 10'b00000_00000;
		Dplus[470] = 10'b00000_00000;
		Dplus[471] = 10'b00000_00000;
		Dplus[472] = 10'b00000_00000;
		Dplus[473] = 10'b00000_00000;
		Dplus[474] = 10'b00000_00000;
		Dplus[475] = 10'b00000_00000;
		Dplus[476] = 10'b00000_00000;
		Dplus[477] = 10'b00000_00000;
		Dplus[478] = 10'b00000_00000;
		Dplus[479] = 10'b00000_00000;
		Dplus[480] = 10'b00000_00000;
		Dplus[481] = 10'b00000_00000;
		Dplus[482] = 10'b00000_00000;
		Dplus[483] = 10'b00000_00000;
		Dplus[484] = 10'b00000_00000;
		Dplus[485] = 10'b00000_00000;
		Dplus[486] = 10'b00000_00000;
		Dplus[487] = 10'b00000_00000;
		Dplus[488] = 10'b00000_00000;
		Dplus[489] = 10'b00000_00000;
		Dplus[490] = 10'b00000_00000;
		Dplus[491] = 10'b00000_00000;
		Dplus[492] = 10'b00000_00000;
		Dplus[493] = 10'b00000_00000;
		Dplus[494] = 10'b00000_00000;
		Dplus[495] = 10'b00000_00000;
		Dplus[496] = 10'b00000_00000;
		Dplus[497] = 10'b00000_00000;
		Dplus[498] = 10'b00000_00000;
		Dplus[499] = 10'b00000_00000;
		Dplus[500] = 10'b00000_00000;
		Dplus[501] = 10'b00000_00000;
		Dplus[502] = 10'b00000_00000;
		Dplus[503] = 10'b00000_00000;
		Dplus[504] = 10'b00000_00000;
		Dplus[505] = 10'b00000_00000;
		Dplus[506] = 10'b00000_00000;
		Dplus[507] = 10'b00000_00000;
		Dplus[508] = 10'b00000_00000;
		Dplus[509] = 10'b00000_00000;
		Dplus[510] = 10'b00000_00000;
		Dplus[511] = 10'b00000_00000;
end
endmodule
