module Tables();
	reg [13:0] Dplus[255:0];
	reg [13:0] Dminus[255:0];
	reg [6:0] DminusInteger[63:0];
	reg [6:0] DplusInteger[63:0];
	initial begin
		Dminus[1] = 14'b1111000_0111100;
		Dminus[2] = 14'b1111001_0111011;
		Dminus[3] = 14'b1111010_0000110;
		Dminus[4] = 14'b1111010_0111010;
		Dminus[5] = 14'b1111010_1100011;
		Dminus[6] = 14'b1111011_0000100;
		Dminus[7] = 14'b1111011_0100000;
		Dminus[8] = 14'b1111011_0111000;
		Dminus[9] = 14'b1111011_1001110;
		Dminus[10] = 14'b1111011_1100001;
		Dminus[11] = 14'b1111011_1110010;
		Dminus[12] = 14'b1111100_0000001;
		Dminus[13] = 14'b1111100_0010000;
		Dminus[14] = 14'b1111100_0011101;
		Dminus[15] = 14'b1111100_0101001;
		Dminus[16] = 14'b1111100_0110100;
		Dminus[17] = 14'b1111100_0111111;
		Dminus[18] = 14'b1111100_1001001;
		Dminus[19] = 14'b1111100_1010011;
		Dminus[20] = 14'b1111100_1011100;
		Dminus[21] = 14'b1111100_1100100;
		Dminus[22] = 14'b1111100_1101100;
		Dminus[23] = 14'b1111100_1110100;
		Dminus[24] = 14'b1111100_1111011;
		Dminus[25] = 14'b1111101_0000010;
		Dminus[26] = 14'b1111101_0001001;
		Dminus[27] = 14'b1111101_0010000;
		Dminus[28] = 14'b1111101_0010110;
		Dminus[29] = 14'b1111101_0011100;
		Dminus[30] = 14'b1111101_0100010;
		Dminus[31] = 14'b1111101_0100111;
		Dminus[32] = 14'b1111101_0101101;
		Dminus[33] = 14'b1111101_0110010;
		Dminus[34] = 14'b1111101_0110111;
		Dminus[35] = 14'b1111101_0111100;
		Dminus[36] = 14'b1111101_1000000;
		Dminus[37] = 14'b1111101_1000101;
		Dminus[38] = 14'b1111101_1001001;
		Dminus[39] = 14'b1111101_1001110;
		Dminus[40] = 14'b1111101_1010010;
		Dminus[41] = 14'b1111101_1010110;
		Dminus[42] = 14'b1111101_1011010;
		Dminus[43] = 14'b1111101_1011110;
		Dminus[44] = 14'b1111101_1100010;
		Dminus[45] = 14'b1111101_1100101;
		Dminus[46] = 14'b1111101_1101001;
		Dminus[47] = 14'b1111101_1101100;
		Dminus[48] = 14'b1111101_1110000;
		Dminus[49] = 14'b1111101_1110011;
		Dminus[50] = 14'b1111101_1110110;
		Dminus[51] = 14'b1111101_1111001;
		Dminus[52] = 14'b1111101_1111101;
		Dminus[53] = 14'b1111110_0000000;
		Dminus[54] = 14'b1111110_0000011;
		Dminus[55] = 14'b1111110_0000110;
		Dminus[56] = 14'b1111110_0001000;
		Dminus[57] = 14'b1111110_0001011;
		Dminus[58] = 14'b1111110_0001110;
		Dminus[59] = 14'b1111110_0010001;
		Dminus[60] = 14'b1111110_0010011;
		Dminus[61] = 14'b1111110_0010110;
		Dminus[62] = 14'b1111110_0011000;
		Dminus[63] = 14'b1111110_0011011;
		Dminus[64] = 14'b1111110_0011101;
		Dminus[65] = 14'b1111110_0100000;
		Dminus[66] = 14'b1111110_0100010;
		Dminus[67] = 14'b1111110_0100100;
		Dminus[68] = 14'b1111110_0100111;
		Dminus[69] = 14'b1111110_0101001;
		Dminus[70] = 14'b1111110_0101011;
		Dminus[71] = 14'b1111110_0101101;
		Dminus[72] = 14'b1111110_0101111;
		Dminus[73] = 14'b1111110_0110001;
		Dminus[74] = 14'b1111110_0110011;
		Dminus[75] = 14'b1111110_0110101;
		Dminus[76] = 14'b1111110_0110111;
		Dminus[77] = 14'b1111110_0111001;
		Dminus[78] = 14'b1111110_0111011;
		Dminus[79] = 14'b1111110_0111101;
		Dminus[80] = 14'b1111110_0111111;
		Dminus[81] = 14'b1111110_1000001;
		Dminus[82] = 14'b1111110_1000011;
		Dminus[83] = 14'b1111110_1000100;
		Dminus[84] = 14'b1111110_1000110;
		Dminus[85] = 14'b1111110_1001000;
		Dminus[86] = 14'b1111110_1001010;
		Dminus[87] = 14'b1111110_1001011;
		Dminus[88] = 14'b1111110_1001101;
		Dminus[89] = 14'b1111110_1001110;
		Dminus[90] = 14'b1111110_1010000;
		Dminus[91] = 14'b1111110_1010010;
		Dminus[92] = 14'b1111110_1010011;
		Dminus[93] = 14'b1111110_1010101;
		Dminus[94] = 14'b1111110_1010110;
		Dminus[95] = 14'b1111110_1011000;
		Dminus[96] = 14'b1111110_1011001;
		Dminus[97] = 14'b1111110_1011011;
		Dminus[98] = 14'b1111110_1011100;
		Dminus[99] = 14'b1111110_1011110;
		Dminus[100] = 14'b1111110_1011111;
		Dminus[101] = 14'b1111110_1100000;
		Dminus[102] = 14'b1111110_1100010;
		Dminus[103] = 14'b1111110_1100011;
		Dminus[104] = 14'b1111110_1100100;
		Dminus[105] = 14'b1111110_1100110;
		Dminus[106] = 14'b1111110_1100111;
		Dminus[107] = 14'b1111110_1101000;
		Dminus[108] = 14'b1111110_1101010;
		Dminus[109] = 14'b1111110_1101011;
		Dminus[110] = 14'b1111110_1101100;
		Dminus[111] = 14'b1111110_1101101;
		Dminus[112] = 14'b1111110_1101110;
		Dminus[113] = 14'b1111110_1110000;
		Dminus[114] = 14'b1111110_1110001;
		Dminus[115] = 14'b1111110_1110010;
		Dminus[116] = 14'b1111110_1110011;
		Dminus[117] = 14'b1111110_1110100;
		Dminus[118] = 14'b1111110_1110101;
		Dminus[119] = 14'b1111110_1110111;
		Dminus[120] = 14'b1111110_1111000;
		Dminus[121] = 14'b1111110_1111001;
		Dminus[122] = 14'b1111110_1111010;
		Dminus[123] = 14'b1111110_1111011;
		Dminus[124] = 14'b1111110_1111100;
		Dminus[125] = 14'b1111110_1111101;
		Dminus[126] = 14'b1111110_1111110;
		Dminus[127] = 14'b1111110_1111111;
		Dminus[128] = 14'b1111111_0000000;
		Dminus[129] = 14'b1111111_0000001;
		Dminus[130] = 14'b1111111_0000010;
		Dminus[131] = 14'b1111111_0000011;
		Dminus[132] = 14'b1111111_0000100;
		Dminus[133] = 14'b1111111_0000101;
		Dminus[134] = 14'b1111111_0000110;
		Dminus[135] = 14'b1111111_0000111;
		Dminus[136] = 14'b1111111_0001000;
		Dminus[137] = 14'b1111111_0001001;
		Dminus[138] = 14'b1111111_0001001;
		Dminus[139] = 14'b1111111_0001010;
		Dminus[140] = 14'b1111111_0001011;
		Dminus[141] = 14'b1111111_0001100;
		Dminus[142] = 14'b1111111_0001101;
		Dminus[143] = 14'b1111111_0001110;
		Dminus[144] = 14'b1111111_0001111;
		Dminus[145] = 14'b1111111_0010000;
		Dminus[146] = 14'b1111111_0010000;
		Dminus[147] = 14'b1111111_0010001;
		Dminus[148] = 14'b1111111_0010010;
		Dminus[149] = 14'b1111111_0010011;
		Dminus[150] = 14'b1111111_0010100;
		Dminus[151] = 14'b1111111_0010100;
		Dminus[152] = 14'b1111111_0010101;
		Dminus[153] = 14'b1111111_0010110;
		Dminus[154] = 14'b1111111_0010111;
		Dminus[155] = 14'b1111111_0011000;
		Dminus[156] = 14'b1111111_0011000;
		Dminus[157] = 14'b1111111_0011001;
		Dminus[158] = 14'b1111111_0011010;
		Dminus[159] = 14'b1111111_0011011;
		Dminus[160] = 14'b1111111_0011011;
		Dminus[161] = 14'b1111111_0011100;
		Dminus[162] = 14'b1111111_0011101;
		Dminus[163] = 14'b1111111_0011101;
		Dminus[164] = 14'b1111111_0011110;
		Dminus[165] = 14'b1111111_0011111;
		Dminus[166] = 14'b1111111_0011111;
		Dminus[167] = 14'b1111111_0100000;
		Dminus[168] = 14'b1111111_0100001;
		Dminus[169] = 14'b1111111_0100010;
		Dminus[170] = 14'b1111111_0100010;
		Dminus[171] = 14'b1111111_0100011;
		Dminus[172] = 14'b1111111_0100100;
		Dminus[173] = 14'b1111111_0100100;
		Dminus[174] = 14'b1111111_0100101;
		Dminus[175] = 14'b1111111_0100101;
		Dminus[176] = 14'b1111111_0100110;
		Dminus[177] = 14'b1111111_0100111;
		Dminus[178] = 14'b1111111_0100111;
		Dminus[179] = 14'b1111111_0101000;
		Dminus[180] = 14'b1111111_0101001;
		Dminus[181] = 14'b1111111_0101001;
		Dminus[182] = 14'b1111111_0101010;
		Dminus[183] = 14'b1111111_0101010;
		Dminus[184] = 14'b1111111_0101011;
		Dminus[185] = 14'b1111111_0101011;
		Dminus[186] = 14'b1111111_0101100;
		Dminus[187] = 14'b1111111_0101101;
		Dminus[188] = 14'b1111111_0101101;
		Dminus[189] = 14'b1111111_0101110;
		Dminus[190] = 14'b1111111_0101110;
		Dminus[191] = 14'b1111111_0101111;
		Dminus[192] = 14'b1111111_0101111;
		Dminus[193] = 14'b1111111_0110000;
		Dminus[194] = 14'b1111111_0110001;
		Dminus[195] = 14'b1111111_0110001;
		Dminus[196] = 14'b1111111_0110010;
		Dminus[197] = 14'b1111111_0110010;
		Dminus[198] = 14'b1111111_0110011;
		Dminus[199] = 14'b1111111_0110011;
		Dminus[200] = 14'b1111111_0110100;
		Dminus[201] = 14'b1111111_0110100;
		Dminus[202] = 14'b1111111_0110101;
		Dminus[203] = 14'b1111111_0110101;
		Dminus[204] = 14'b1111111_0110110;
		Dminus[205] = 14'b1111111_0110110;
		Dminus[206] = 14'b1111111_0110111;
		Dminus[207] = 14'b1111111_0110111;
		Dminus[208] = 14'b1111111_0111000;
		Dminus[209] = 14'b1111111_0111000;
		Dminus[210] = 14'b1111111_0111001;
		Dminus[211] = 14'b1111111_0111001;
		Dminus[212] = 14'b1111111_0111010;
		Dminus[213] = 14'b1111111_0111010;
		Dminus[214] = 14'b1111111_0111010;
		Dminus[215] = 14'b1111111_0111011;
		Dminus[216] = 14'b1111111_0111011;
		Dminus[217] = 14'b1111111_0111100;
		Dminus[218] = 14'b1111111_0111100;
		Dminus[219] = 14'b1111111_0111101;
		Dminus[220] = 14'b1111111_0111101;
		Dminus[221] = 14'b1111111_0111110;
		Dminus[222] = 14'b1111111_0111110;
		Dminus[223] = 14'b1111111_0111110;
		Dminus[224] = 14'b1111111_0111111;
		Dminus[225] = 14'b1111111_0111111;
		Dminus[226] = 14'b1111111_1000000;
		Dminus[227] = 14'b1111111_1000000;
		Dminus[228] = 14'b1111111_1000001;
		Dminus[229] = 14'b1111111_1000001;
		Dminus[230] = 14'b1111111_1000001;
		Dminus[231] = 14'b1111111_1000010;
		Dminus[232] = 14'b1111111_1000010;
		Dminus[233] = 14'b1111111_1000011;
		Dminus[234] = 14'b1111111_1000011;
		Dminus[235] = 14'b1111111_1000011;
		Dminus[236] = 14'b1111111_1000100;
		Dminus[237] = 14'b1111111_1000100;
		Dminus[238] = 14'b1111111_1000100;
		Dminus[239] = 14'b1111111_1000101;
		Dminus[240] = 14'b1111111_1000101;
		Dminus[241] = 14'b1111111_1000110;
		Dminus[242] = 14'b1111111_1000110;
		Dminus[243] = 14'b1111111_1000110;
		Dminus[244] = 14'b1111111_1000111;
		Dminus[245] = 14'b1111111_1000111;
		Dminus[246] = 14'b1111111_1000111;
		Dminus[247] = 14'b1111111_1001000;
		Dminus[248] = 14'b1111111_1001000;
		Dminus[249] = 14'b1111111_1001000;
		Dminus[250] = 14'b1111111_1001001;
		Dminus[251] = 14'b1111111_1001001;
		Dminus[252] = 14'b1111111_1001010;
		Dminus[253] = 14'b1111111_1001010;
		Dminus[254] = 14'b1111111_1001010;
		Dminus[255] = 14'b1111111_1001011;
		Dplus[1] = 14'b0000001_0000000;
		Dplus[2] = 14'b0000000_1111111;
		Dplus[3] = 14'b0000000_1111111;
		Dplus[4] = 14'b0000000_1111110;
		Dplus[5] = 14'b0000000_1111110;
		Dplus[6] = 14'b0000000_1111101;
		Dplus[7] = 14'b0000000_1111101;
		Dplus[8] = 14'b0000000_1111100;
		Dplus[9] = 14'b0000000_1111100;
		Dplus[10] = 14'b0000000_1111011;
		Dplus[11] = 14'b0000000_1111011;
		Dplus[12] = 14'b0000000_1111010;
		Dplus[13] = 14'b0000000_1111010;
		Dplus[14] = 14'b0000000_1111001;
		Dplus[15] = 14'b0000000_1111001;
		Dplus[16] = 14'b0000000_1111000;
		Dplus[17] = 14'b0000000_1111000;
		Dplus[18] = 14'b0000000_1110111;
		Dplus[19] = 14'b0000000_1110111;
		Dplus[20] = 14'b0000000_1110110;
		Dplus[21] = 14'b0000000_1110110;
		Dplus[22] = 14'b0000000_1110101;
		Dplus[23] = 14'b0000000_1110101;
		Dplus[24] = 14'b0000000_1110100;
		Dplus[25] = 14'b0000000_1110100;
		Dplus[26] = 14'b0000000_1110011;
		Dplus[27] = 14'b0000000_1110011;
		Dplus[28] = 14'b0000000_1110011;
		Dplus[29] = 14'b0000000_1110010;
		Dplus[30] = 14'b0000000_1110010;
		Dplus[31] = 14'b0000000_1110001;
		Dplus[32] = 14'b0000000_1110001;
		Dplus[33] = 14'b0000000_1110000;
		Dplus[34] = 14'b0000000_1110000;
		Dplus[35] = 14'b0000000_1101111;
		Dplus[36] = 14'b0000000_1101111;
		Dplus[37] = 14'b0000000_1101110;
		Dplus[38] = 14'b0000000_1101110;
		Dplus[39] = 14'b0000000_1101110;
		Dplus[40] = 14'b0000000_1101101;
		Dplus[41] = 14'b0000000_1101101;
		Dplus[42] = 14'b0000000_1101100;
		Dplus[43] = 14'b0000000_1101100;
		Dplus[44] = 14'b0000000_1101011;
		Dplus[45] = 14'b0000000_1101011;
		Dplus[46] = 14'b0000000_1101010;
		Dplus[47] = 14'b0000000_1101010;
		Dplus[48] = 14'b0000000_1101010;
		Dplus[49] = 14'b0000000_1101001;
		Dplus[50] = 14'b0000000_1101001;
		Dplus[51] = 14'b0000000_1101000;
		Dplus[52] = 14'b0000000_1101000;
		Dplus[53] = 14'b0000000_1100111;
		Dplus[54] = 14'b0000000_1100111;
		Dplus[55] = 14'b0000000_1100111;
		Dplus[56] = 14'b0000000_1100110;
		Dplus[57] = 14'b0000000_1100110;
		Dplus[58] = 14'b0000000_1100101;
		Dplus[59] = 14'b0000000_1100101;
		Dplus[60] = 14'b0000000_1100100;
		Dplus[61] = 14'b0000000_1100100;
		Dplus[62] = 14'b0000000_1100100;
		Dplus[63] = 14'b0000000_1100011;
		Dplus[64] = 14'b0000000_1100011;
		Dplus[65] = 14'b0000000_1100010;
		Dplus[66] = 14'b0000000_1100010;
		Dplus[67] = 14'b0000000_1100010;
		Dplus[68] = 14'b0000000_1100001;
		Dplus[69] = 14'b0000000_1100001;
		Dplus[70] = 14'b0000000_1100000;
		Dplus[71] = 14'b0000000_1100000;
		Dplus[72] = 14'b0000000_1011111;
		Dplus[73] = 14'b0000000_1011111;
		Dplus[74] = 14'b0000000_1011111;
		Dplus[75] = 14'b0000000_1011110;
		Dplus[76] = 14'b0000000_1011110;
		Dplus[77] = 14'b0000000_1011101;
		Dplus[78] = 14'b0000000_1011101;
		Dplus[79] = 14'b0000000_1011101;
		Dplus[80] = 14'b0000000_1011100;
		Dplus[81] = 14'b0000000_1011100;
		Dplus[82] = 14'b0000000_1011100;
		Dplus[83] = 14'b0000000_1011011;
		Dplus[84] = 14'b0000000_1011011;
		Dplus[85] = 14'b0000000_1011010;
		Dplus[86] = 14'b0000000_1011010;
		Dplus[87] = 14'b0000000_1011010;
		Dplus[88] = 14'b0000000_1011001;
		Dplus[89] = 14'b0000000_1011001;
		Dplus[90] = 14'b0000000_1011000;
		Dplus[91] = 14'b0000000_1011000;
		Dplus[92] = 14'b0000000_1011000;
		Dplus[93] = 14'b0000000_1010111;
		Dplus[94] = 14'b0000000_1010111;
		Dplus[95] = 14'b0000000_1010111;
		Dplus[96] = 14'b0000000_1010110;
		Dplus[97] = 14'b0000000_1010110;
		Dplus[98] = 14'b0000000_1010101;
		Dplus[99] = 14'b0000000_1010101;
		Dplus[100] = 14'b0000000_1010101;
		Dplus[101] = 14'b0000000_1010100;
		Dplus[102] = 14'b0000000_1010100;
		Dplus[103] = 14'b0000000_1010100;
		Dplus[104] = 14'b0000000_1010011;
		Dplus[105] = 14'b0000000_1010011;
		Dplus[106] = 14'b0000000_1010011;
		Dplus[107] = 14'b0000000_1010010;
		Dplus[108] = 14'b0000000_1010010;
		Dplus[109] = 14'b0000000_1010001;
		Dplus[110] = 14'b0000000_1010001;
		Dplus[111] = 14'b0000000_1010001;
		Dplus[112] = 14'b0000000_1010000;
		Dplus[113] = 14'b0000000_1010000;
		Dplus[114] = 14'b0000000_1010000;
		Dplus[115] = 14'b0000000_1001111;
		Dplus[116] = 14'b0000000_1001111;
		Dplus[117] = 14'b0000000_1001111;
		Dplus[118] = 14'b0000000_1001110;
		Dplus[119] = 14'b0000000_1001110;
		Dplus[120] = 14'b0000000_1001110;
		Dplus[121] = 14'b0000000_1001101;
		Dplus[122] = 14'b0000000_1001101;
		Dplus[123] = 14'b0000000_1001101;
		Dplus[124] = 14'b0000000_1001100;
		Dplus[125] = 14'b0000000_1001100;
		Dplus[126] = 14'b0000000_1001100;
		Dplus[127] = 14'b0000000_1001011;
		Dplus[128] = 14'b0000000_1001011;
		Dplus[129] = 14'b0000000_1001011;
		Dplus[130] = 14'b0000000_1001010;
		Dplus[131] = 14'b0000000_1001010;
		Dplus[132] = 14'b0000000_1001010;
		Dplus[133] = 14'b0000000_1001001;
		Dplus[134] = 14'b0000000_1001001;
		Dplus[135] = 14'b0000000_1001001;
		Dplus[136] = 14'b0000000_1001000;
		Dplus[137] = 14'b0000000_1001000;
		Dplus[138] = 14'b0000000_1001000;
		Dplus[139] = 14'b0000000_1000111;
		Dplus[140] = 14'b0000000_1000111;
		Dplus[141] = 14'b0000000_1000111;
		Dplus[142] = 14'b0000000_1000110;
		Dplus[143] = 14'b0000000_1000110;
		Dplus[144] = 14'b0000000_1000110;
		Dplus[145] = 14'b0000000_1000101;
		Dplus[146] = 14'b0000000_1000101;
		Dplus[147] = 14'b0000000_1000101;
		Dplus[148] = 14'b0000000_1000100;
		Dplus[149] = 14'b0000000_1000100;
		Dplus[150] = 14'b0000000_1000100;
		Dplus[151] = 14'b0000000_1000100;
		Dplus[152] = 14'b0000000_1000011;
		Dplus[153] = 14'b0000000_1000011;
		Dplus[154] = 14'b0000000_1000011;
		Dplus[155] = 14'b0000000_1000010;
		Dplus[156] = 14'b0000000_1000010;
		Dplus[157] = 14'b0000000_1000010;
		Dplus[158] = 14'b0000000_1000001;
		Dplus[159] = 14'b0000000_1000001;
		Dplus[160] = 14'b0000000_1000001;
		Dplus[161] = 14'b0000000_1000001;
		Dplus[162] = 14'b0000000_1000000;
		Dplus[163] = 14'b0000000_1000000;
		Dplus[164] = 14'b0000000_1000000;
		Dplus[165] = 14'b0000000_0111111;
		Dplus[166] = 14'b0000000_0111111;
		Dplus[167] = 14'b0000000_0111111;
		Dplus[168] = 14'b0000000_0111110;
		Dplus[169] = 14'b0000000_0111110;
		Dplus[170] = 14'b0000000_0111110;
		Dplus[171] = 14'b0000000_0111110;
		Dplus[172] = 14'b0000000_0111101;
		Dplus[173] = 14'b0000000_0111101;
		Dplus[174] = 14'b0000000_0111101;
		Dplus[175] = 14'b0000000_0111100;
		Dplus[176] = 14'b0000000_0111100;
		Dplus[177] = 14'b0000000_0111100;
		Dplus[178] = 14'b0000000_0111100;
		Dplus[179] = 14'b0000000_0111011;
		Dplus[180] = 14'b0000000_0111011;
		Dplus[181] = 14'b0000000_0111011;
		Dplus[182] = 14'b0000000_0111011;
		Dplus[183] = 14'b0000000_0111010;
		Dplus[184] = 14'b0000000_0111010;
		Dplus[185] = 14'b0000000_0111010;
		Dplus[186] = 14'b0000000_0111001;
		Dplus[187] = 14'b0000000_0111001;
		Dplus[188] = 14'b0000000_0111001;
		Dplus[189] = 14'b0000000_0111001;
		Dplus[190] = 14'b0000000_0111000;
		Dplus[191] = 14'b0000000_0111000;
		Dplus[192] = 14'b0000000_0111000;
		Dplus[193] = 14'b0000000_0111000;
		Dplus[194] = 14'b0000000_0110111;
		Dplus[195] = 14'b0000000_0110111;
		Dplus[196] = 14'b0000000_0110111;
		Dplus[197] = 14'b0000000_0110111;
		Dplus[198] = 14'b0000000_0110110;
		Dplus[199] = 14'b0000000_0110110;
		Dplus[200] = 14'b0000000_0110110;
		Dplus[201] = 14'b0000000_0110110;
		Dplus[202] = 14'b0000000_0110101;
		Dplus[203] = 14'b0000000_0110101;
		Dplus[204] = 14'b0000000_0110101;
		Dplus[205] = 14'b0000000_0110101;
		Dplus[206] = 14'b0000000_0110100;
		Dplus[207] = 14'b0000000_0110100;
		Dplus[208] = 14'b0000000_0110100;
		Dplus[209] = 14'b0000000_0110100;
		Dplus[210] = 14'b0000000_0110011;
		Dplus[211] = 14'b0000000_0110011;
		Dplus[212] = 14'b0000000_0110011;
		Dplus[213] = 14'b0000000_0110011;
		Dplus[214] = 14'b0000000_0110010;
		Dplus[215] = 14'b0000000_0110010;
		Dplus[216] = 14'b0000000_0110010;
		Dplus[217] = 14'b0000000_0110010;
		Dplus[218] = 14'b0000000_0110001;
		Dplus[219] = 14'b0000000_0110001;
		Dplus[220] = 14'b0000000_0110001;
		Dplus[221] = 14'b0000000_0110001;
		Dplus[222] = 14'b0000000_0110001;
		Dplus[223] = 14'b0000000_0110000;
		Dplus[224] = 14'b0000000_0110000;
		Dplus[225] = 14'b0000000_0110000;
		Dplus[226] = 14'b0000000_0110000;
		Dplus[227] = 14'b0000000_0101111;
		Dplus[228] = 14'b0000000_0101111;
		Dplus[229] = 14'b0000000_0101111;
		Dplus[230] = 14'b0000000_0101111;
		Dplus[231] = 14'b0000000_0101110;
		Dplus[232] = 14'b0000000_0101110;
		Dplus[233] = 14'b0000000_0101110;
		Dplus[234] = 14'b0000000_0101110;
		Dplus[235] = 14'b0000000_0101110;
		Dplus[236] = 14'b0000000_0101101;
		Dplus[237] = 14'b0000000_0101101;
		Dplus[238] = 14'b0000000_0101101;
		Dplus[239] = 14'b0000000_0101101;
		Dplus[240] = 14'b0000000_0101101;
		Dplus[241] = 14'b0000000_0101100;
		Dplus[242] = 14'b0000000_0101100;
		Dplus[243] = 14'b0000000_0101100;
		Dplus[244] = 14'b0000000_0101100;
		Dplus[245] = 14'b0000000_0101011;
		Dplus[246] = 14'b0000000_0101011;
		Dplus[247] = 14'b0000000_0101011;
		Dplus[248] = 14'b0000000_0101011;
		Dplus[249] = 14'b0000000_0101011;
		Dplus[250] = 14'b0000000_0101010;
		Dplus[251] = 14'b0000000_0101010;
		Dplus[252] = 14'b0000000_0101010;
		Dplus[253] = 14'b0000000_0101010;
		Dplus[254] = 14'b0000000_0101010;
		Dplus[255] = 14'b0000000_0101001;
		DplusInteger[2] = 14'b0000000_0101001;
		DplusInteger[3] = 14'b0000000_0010110;
		DplusInteger[4] = 14'b0000000_0001011;
		DplusInteger[5] = 14'b0000000_0000110;
		DplusInteger[6] = 14'b0000000_0000011;
		DplusInteger[7] = 14'b0000000_0000001;
		DplusInteger[8] = 14'b0000000_0000001;
		DplusInteger[9] = 14'b0000000_0000000;
		DplusInteger[10] = 14'b0000000_0000000;
		DplusInteger[11] = 14'b0000000_0000000;
		DplusInteger[12] = 14'b0000000_0000000;
		DplusInteger[13] = 14'b0000000_0000000;
		DplusInteger[14] = 14'b0000000_0000000;
		DplusInteger[15] = 14'b0000000_0000000;
		DplusInteger[16] = 14'b0000000_0000000;
		DplusInteger[17] = 14'b0000000_0000000;
		DplusInteger[18] = 14'b0000000_0000000;
		DplusInteger[19] = 14'b0000000_0000000;
		DplusInteger[20] = 14'b0000000_0000000;
		DplusInteger[21] = 14'b0000000_0000000;
		DplusInteger[22] = 14'b0000000_0000000;
		DplusInteger[23] = 14'b0000000_0000000;
		DplusInteger[24] = 14'b0000000_0000000;
		DplusInteger[25] = 14'b0000000_0000000;
		DplusInteger[26] = 14'b0000000_0000000;
		DplusInteger[27] = 14'b0000000_0000000;
		DplusInteger[28] = 14'b0000000_0000000;
		DplusInteger[29] = 14'b0000000_0000000;
		DplusInteger[30] = 14'b0000000_0000000;
		DplusInteger[31] = 14'b0000000_0000000;
		DplusInteger[32] = 14'b0000000_0000000;
		DplusInteger[33] = 14'b0000000_0000000;
		DplusInteger[34] = 14'b0000000_0000000;
		DplusInteger[35] = 14'b0000000_0000000;
		DplusInteger[36] = 14'b0000000_0000000;
		DplusInteger[37] = 14'b0000000_0000000;
		DplusInteger[38] = 14'b0000000_0000000;
		DplusInteger[39] = 14'b0000000_0000000;
		DplusInteger[40] = 14'b0000000_0000000;
		DplusInteger[41] = 14'b0000000_0000000;
		DplusInteger[42] = 14'b0000000_0000000;
		DplusInteger[43] = 14'b0000000_0000000;
		DplusInteger[44] = 14'b0000000_0000000;
		DplusInteger[45] = 14'b0000000_0000000;
		DplusInteger[46] = 14'b0000000_0000000;
		DplusInteger[47] = 14'b0000000_0000000;
		DplusInteger[48] = 14'b0000000_0000000;
		DplusInteger[49] = 14'b0000000_0000000;
		DplusInteger[50] = 14'b0000000_0000000;
		DplusInteger[51] = 14'b0000000_0000000;
		DplusInteger[52] = 14'b0000000_0000000;
		DplusInteger[53] = 14'b0000000_0000000;
		DplusInteger[54] = 14'b0000000_0000000;
		DplusInteger[55] = 14'b0000000_0000000;
		DplusInteger[56] = 14'b0000000_0000000;
		DplusInteger[57] = 14'b0000000_0000000;
		DplusInteger[58] = 14'b0000000_0000000;
		DplusInteger[59] = 14'b0000000_0000000;
		DplusInteger[60] = 14'b0000000_0000000;
		DplusInteger[61] = 14'b0000000_0000000;
		DplusInteger[62] = 14'b0000000_0000000;
		DplusInteger[63] = 14'b0000000_0000000;
		DminusInteger[2] = 14'b1111111_1001011;
		DminusInteger[3] = 14'b1111111_1100111;
		DminusInteger[4] = 14'b1111111_1110100;
		DminusInteger[5] = 14'b1111111_1111010;
		DminusInteger[6] = 14'b1111111_1111101;
		DminusInteger[7] = 14'b1111111_1111111;
		DminusInteger[8] = 14'b1111111_1111111;
		DminusInteger[9] = 14'b0000000_0000000;
		DminusInteger[10] = 14'b0000000_0000000;
		DminusInteger[11] = 14'b0000000_0000000;
		DminusInteger[12] = 14'b0000000_0000000;
		DminusInteger[13] = 14'b0000000_0000000;
		DminusInteger[14] = 14'b0000000_0000000;
		DminusInteger[15] = 14'b0000000_0000000;
		DminusInteger[16] = 14'b0000000_0000000;
		DminusInteger[17] = 14'b0000000_0000000;
		DminusInteger[18] = 14'b0000000_0000000;
		DminusInteger[19] = 14'b0000000_0000000;
		DminusInteger[20] = 14'b0000000_0000000;
		DminusInteger[21] = 14'b0000000_0000000;
		DminusInteger[22] = 14'b0000000_0000000;
		DminusInteger[23] = 14'b0000000_0000000;
		DminusInteger[24] = 14'b0000000_0000000;
		DminusInteger[25] = 14'b0000000_0000000;
		DminusInteger[26] = 14'b0000000_0000000;
		DminusInteger[27] = 14'b0000000_0000000;
		DminusInteger[28] = 14'b0000000_0000000;
		DminusInteger[29] = 14'b0000000_0000000;
		DminusInteger[30] = 14'b0000000_0000000;
		DminusInteger[31] = 14'b0000000_0000000;
		DminusInteger[32] = 14'b0000000_0000000;
		DminusInteger[33] = 14'b0000000_0000000;
		DminusInteger[34] = 14'b0000000_0000000;
		DminusInteger[35] = 14'b0000000_0000000;
		DminusInteger[36] = 14'b0000000_0000000;
		DminusInteger[37] = 14'b0000000_0000000;
		DminusInteger[38] = 14'b0000000_0000000;
		DminusInteger[39] = 14'b0000000_0000000;
		DminusInteger[40] = 14'b0000000_0000000;
		DminusInteger[41] = 14'b0000000_0000000;
		DminusInteger[42] = 14'b0000000_0000000;
		DminusInteger[43] = 14'b0000000_0000000;
		DminusInteger[44] = 14'b0000000_0000000;
		DminusInteger[45] = 14'b0000000_0000000;
		DminusInteger[46] = 14'b0000000_0000000;
		DminusInteger[47] = 14'b0000000_0000000;
		DminusInteger[48] = 14'b0000000_0000000;
		DminusInteger[49] = 14'b0000000_0000000;
		DminusInteger[50] = 14'b0000000_0000000;
		DminusInteger[51] = 14'b0000000_0000000;
		DminusInteger[52] = 14'b0000000_0000000;
		DminusInteger[53] = 14'b0000000_0000000;
		DminusInteger[54] = 14'b0000000_0000000;
		DminusInteger[55] = 14'b0000000_0000000;
		DminusInteger[56] = 14'b0000000_0000000;
		DminusInteger[57] = 14'b0000000_0000000;
		DminusInteger[58] = 14'b0000000_0000000;
		DminusInteger[59] = 14'b0000000_0000000;
		DminusInteger[60] = 14'b0000000_0000000;
		DminusInteger[61] = 14'b0000000_0000000;
		DminusInteger[62] = 14'b0000000_0000000;
		DminusInteger[63] = 14'b0000000_0000000;
end
endmodule
