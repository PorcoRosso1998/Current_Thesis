module Tables();
	reg [7:0] Dplus[31:0];
	reg [7:0] Dminus[31:0];
	reg [3:0] DminusInteger[7:0];
	reg [3:0] DplusInteger[7:0];
	initial begin
		Dminus[1] = 8'b1011_0111;
		Dminus[2] = 8'b1100_0111;
		Dminus[3] = 8'b1100_1111;
		Dminus[4] = 8'b1101_0110;
		Dminus[5] = 8'b1101_1010;
		Dminus[6] = 8'b1101_1110;
		Dminus[7] = 8'b1110_0001;
		Dminus[8] = 8'b1110_0100;
		Dminus[9] = 8'b1110_0110;
		Dminus[10] = 8'b1110_1000;
		Dminus[11] = 8'b1110_1010;
		Dminus[12] = 8'b1110_1011;
		Dminus[13] = 8'b1110_1101;
		Dminus[14] = 8'b1110_1110;
		Dminus[15] = 8'b1110_1111;
		Dminus[16] = 8'b1111_0000;
		Dminus[17] = 8'b1111_0001;
		Dminus[18] = 8'b1111_0010;
		Dminus[19] = 8'b1111_0011;
		Dminus[20] = 8'b1111_0011;
		Dminus[21] = 8'b1111_0100;
		Dminus[22] = 8'b1111_0101;
		Dminus[23] = 8'b1111_0101;
		Dminus[24] = 8'b1111_0110;
		Dminus[25] = 8'b1111_0110;
		Dminus[26] = 8'b1111_0111;
		Dminus[27] = 8'b1111_0111;
		Dminus[28] = 8'b1111_1000;
		Dminus[29] = 8'b1111_1000;
		Dminus[30] = 8'b1111_1001;
		Dminus[31] = 8'b1111_1001;
		Dplus[1] = 8'b0001_0000;
		Dplus[2] = 8'b0000_1111;
		Dplus[3] = 8'b0000_1111;
		Dplus[4] = 8'b0000_1110;
		Dplus[5] = 8'b0000_1110;
		Dplus[6] = 8'b0000_1101;
		Dplus[7] = 8'b0000_1101;
		Dplus[8] = 8'b0000_1100;
		Dplus[9] = 8'b0000_1100;
		Dplus[10] = 8'b0000_1100;
		Dplus[11] = 8'b0000_1011;
		Dplus[12] = 8'b0000_1011;
		Dplus[13] = 8'b0000_1010;
		Dplus[14] = 8'b0000_1010;
		Dplus[15] = 8'b0000_1010;
		Dplus[16] = 8'b0000_1001;
		Dplus[17] = 8'b0000_1001;
		Dplus[18] = 8'b0000_1001;
		Dplus[19] = 8'b0000_1000;
		Dplus[20] = 8'b0000_1000;
		Dplus[21] = 8'b0000_1000;
		Dplus[22] = 8'b0000_1000;
		Dplus[23] = 8'b0000_0111;
		Dplus[24] = 8'b0000_0111;
		Dplus[25] = 8'b0000_0111;
		Dplus[26] = 8'b0000_0110;
		Dplus[27] = 8'b0000_0110;
		Dplus[28] = 8'b0000_0110;
		Dplus[29] = 8'b0000_0110;
		Dplus[30] = 8'b0000_0110;
		Dplus[31] = 8'b0000_0101;
		DplusInteger[2] = 8'b0000_0101;
		DplusInteger[3] = 8'b0000_0011;
		DplusInteger[4] = 8'b0000_0001;
		DplusInteger[5] = 8'b0000_0001;
		DplusInteger[6] = 8'b0000_0000;
		DplusInteger[7] = 8'b0000_0000;
		DminusInteger[2] = 8'b1111_1001;
		DminusInteger[3] = 8'b1111_1101;
		DminusInteger[4] = 8'b1111_1111;
		DminusInteger[5] = 8'b1111_1111;
		DminusInteger[6] = 8'b0000_0000;
		DminusInteger[7] = 8'b0000_0000;
end
endmodule
