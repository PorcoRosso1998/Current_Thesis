module Tables();
	reg [7:0] logarithm_table[127:0];
	reg [7:0] Dplus[127:0];
	reg [7:0] Dminus[127:0];
	initial begin
		logarithm_table[1] = 8'b1100_0000;
		logarithm_table[2] = 8'b1101_0000;
		logarithm_table[3] = 8'b1101_1001;
		logarithm_table[4] = 8'b1110_0000;
		logarithm_table[5] = 8'b1110_0101;
		logarithm_table[6] = 8'b1110_1001;
		logarithm_table[7] = 8'b1110_1101;
		logarithm_table[8] = 8'b1111_0000;
		logarithm_table[9] = 8'b1111_0011;
		logarithm_table[10] = 8'b1111_0101;
		logarithm_table[11] = 8'b1111_0111;
		logarithm_table[12] = 8'b1111_1001;
		logarithm_table[13] = 8'b1111_1011;
		logarithm_table[14] = 8'b1111_1101;
		logarithm_table[15] = 8'b1111_1111;
		logarithm_table[16] = 8'b0000_0000;
		logarithm_table[17] = 8'b0000_0001;
		logarithm_table[18] = 8'b0000_0011;
		logarithm_table[19] = 8'b0000_0100;
		logarithm_table[20] = 8'b0000_0101;
		logarithm_table[21] = 8'b0000_0110;
		logarithm_table[22] = 8'b0000_0111;
		logarithm_table[23] = 8'b0000_1000;
		logarithm_table[24] = 8'b0000_1001;
		logarithm_table[25] = 8'b0000_1010;
		logarithm_table[26] = 8'b0000_1011;
		logarithm_table[27] = 8'b0000_1100;
		logarithm_table[28] = 8'b0000_1101;
		logarithm_table[29] = 8'b0000_1110;
		logarithm_table[30] = 8'b0000_1111;
		logarithm_table[31] = 8'b0000_1111;
		logarithm_table[32] = 8'b0001_0000;
		logarithm_table[33] = 8'b0001_0001;
		logarithm_table[34] = 8'b0001_0001;
		logarithm_table[35] = 8'b0001_0010;
		logarithm_table[36] = 8'b0001_0011;
		logarithm_table[37] = 8'b0001_0011;
		logarithm_table[38] = 8'b0001_0100;
		logarithm_table[39] = 8'b0001_0101;
		logarithm_table[40] = 8'b0001_0101;
		logarithm_table[41] = 8'b0001_0110;
		logarithm_table[42] = 8'b0001_0110;
		logarithm_table[43] = 8'b0001_0111;
		logarithm_table[44] = 8'b0001_0111;
		logarithm_table[45] = 8'b0001_1000;
		logarithm_table[46] = 8'b0001_1000;
		logarithm_table[47] = 8'b0001_1001;
		logarithm_table[48] = 8'b0001_1001;
		logarithm_table[49] = 8'b0001_1010;
		logarithm_table[50] = 8'b0001_1010;
		logarithm_table[51] = 8'b0001_1011;
		logarithm_table[52] = 8'b0001_1011;
		logarithm_table[53] = 8'b0001_1100;
		logarithm_table[54] = 8'b0001_1100;
		logarithm_table[55] = 8'b0001_1101;
		logarithm_table[56] = 8'b0001_1101;
		logarithm_table[57] = 8'b0001_1101;
		logarithm_table[58] = 8'b0001_1110;
		logarithm_table[59] = 8'b0001_1110;
		logarithm_table[60] = 8'b0001_1111;
		logarithm_table[61] = 8'b0001_1111;
		logarithm_table[62] = 8'b0001_1111;
		logarithm_table[63] = 8'b0010_0000;
		logarithm_table[64] = 8'b0010_0000;
		logarithm_table[65] = 8'b0010_0000;
		logarithm_table[66] = 8'b0010_0001;
		logarithm_table[67] = 8'b0010_0001;
		logarithm_table[68] = 8'b0010_0001;
		logarithm_table[69] = 8'b0010_0010;
		logarithm_table[70] = 8'b0010_0010;
		logarithm_table[71] = 8'b0010_0010;
		logarithm_table[72] = 8'b0010_0011;
		logarithm_table[73] = 8'b0010_0011;
		logarithm_table[74] = 8'b0010_0011;
		logarithm_table[75] = 8'b0010_0100;
		logarithm_table[76] = 8'b0010_0100;
		logarithm_table[77] = 8'b0010_0100;
		logarithm_table[78] = 8'b0010_0101;
		logarithm_table[79] = 8'b0010_0101;
		logarithm_table[80] = 8'b0010_0101;
		logarithm_table[81] = 8'b0010_0101;
		logarithm_table[82] = 8'b0010_0110;
		logarithm_table[83] = 8'b0010_0110;
		logarithm_table[84] = 8'b0010_0110;
		logarithm_table[85] = 8'b0010_0111;
		logarithm_table[86] = 8'b0010_0111;
		logarithm_table[87] = 8'b0010_0111;
		logarithm_table[88] = 8'b0010_0111;
		logarithm_table[89] = 8'b0010_1000;
		logarithm_table[90] = 8'b0010_1000;
		logarithm_table[91] = 8'b0010_1000;
		logarithm_table[92] = 8'b0010_1000;
		logarithm_table[93] = 8'b0010_1001;
		logarithm_table[94] = 8'b0010_1001;
		logarithm_table[95] = 8'b0010_1001;
		logarithm_table[96] = 8'b0010_1001;
		logarithm_table[97] = 8'b0010_1010;
		logarithm_table[98] = 8'b0010_1010;
		logarithm_table[99] = 8'b0010_1010;
		logarithm_table[100] = 8'b0010_1010;
		logarithm_table[101] = 8'b0010_1011;
		logarithm_table[102] = 8'b0010_1011;
		logarithm_table[103] = 8'b0010_1011;
		logarithm_table[104] = 8'b0010_1011;
		logarithm_table[105] = 8'b0010_1011;
		logarithm_table[106] = 8'b0010_1100;
		logarithm_table[107] = 8'b0010_1100;
		logarithm_table[108] = 8'b0010_1100;
		logarithm_table[109] = 8'b0010_1100;
		logarithm_table[110] = 8'b0010_1101;
		logarithm_table[111] = 8'b0010_1101;
		logarithm_table[112] = 8'b0010_1101;
		logarithm_table[113] = 8'b0010_1101;
		logarithm_table[114] = 8'b0010_1101;
		logarithm_table[115] = 8'b0010_1110;
		logarithm_table[116] = 8'b0010_1110;
		logarithm_table[117] = 8'b0010_1110;
		logarithm_table[118] = 8'b0010_1110;
		logarithm_table[119] = 8'b0010_1110;
		logarithm_table[120] = 8'b0010_1111;
		logarithm_table[121] = 8'b0010_1111;
		logarithm_table[122] = 8'b0010_1111;
		logarithm_table[123] = 8'b0010_1111;
		logarithm_table[124] = 8'b0010_1111;
		logarithm_table[125] = 8'b0010_1111;
		logarithm_table[126] = 8'b0011_0000;
		logarithm_table[127] = 8'b0011_0000;
		Dminus[1] = 8'b1011_0111;
		Dminus[2] = 8'b1100_0111;
		Dminus[3] = 8'b1100_1111;
		Dminus[4] = 8'b1101_0110;
		Dminus[5] = 8'b1101_1010;
		Dminus[6] = 8'b1101_1110;
		Dminus[7] = 8'b1110_0001;
		Dminus[8] = 8'b1110_0100;
		Dminus[9] = 8'b1110_0110;
		Dminus[10] = 8'b1110_1000;
		Dminus[11] = 8'b1110_1010;
		Dminus[12] = 8'b1110_1011;
		Dminus[13] = 8'b1110_1101;
		Dminus[14] = 8'b1110_1110;
		Dminus[15] = 8'b1110_1111;
		Dminus[16] = 8'b1111_0000;
		Dminus[17] = 8'b1111_0001;
		Dminus[18] = 8'b1111_0010;
		Dminus[19] = 8'b1111_0011;
		Dminus[20] = 8'b1111_0011;
		Dminus[21] = 8'b1111_0100;
		Dminus[22] = 8'b1111_0101;
		Dminus[23] = 8'b1111_0101;
		Dminus[24] = 8'b1111_0110;
		Dminus[25] = 8'b1111_0110;
		Dminus[26] = 8'b1111_0111;
		Dminus[27] = 8'b1111_0111;
		Dminus[28] = 8'b1111_1000;
		Dminus[29] = 8'b1111_1000;
		Dminus[30] = 8'b1111_1001;
		Dminus[31] = 8'b1111_1001;
		Dminus[32] = 8'b1111_1001;
		Dminus[33] = 8'b1111_1010;
		Dminus[34] = 8'b1111_1010;
		Dminus[35] = 8'b1111_1010;
		Dminus[36] = 8'b1111_1011;
		Dminus[37] = 8'b1111_1011;
		Dminus[38] = 8'b1111_1011;
		Dminus[39] = 8'b1111_1011;
		Dminus[40] = 8'b1111_1100;
		Dminus[41] = 8'b1111_1100;
		Dminus[42] = 8'b1111_1100;
		Dminus[43] = 8'b1111_1100;
		Dminus[44] = 8'b1111_1100;
		Dminus[45] = 8'b1111_1100;
		Dminus[46] = 8'b1111_1101;
		Dminus[47] = 8'b1111_1101;
		Dminus[48] = 8'b1111_1101;
		Dminus[49] = 8'b1111_1101;
		Dminus[50] = 8'b1111_1101;
		Dminus[51] = 8'b1111_1101;
		Dminus[52] = 8'b1111_1101;
		Dminus[53] = 8'b1111_1110;
		Dminus[54] = 8'b1111_1110;
		Dminus[55] = 8'b1111_1110;
		Dminus[56] = 8'b1111_1110;
		Dminus[57] = 8'b1111_1110;
		Dminus[58] = 8'b1111_1110;
		Dminus[59] = 8'b1111_1110;
		Dminus[60] = 8'b1111_1110;
		Dminus[61] = 8'b1111_1110;
		Dminus[62] = 8'b1111_1110;
		Dminus[63] = 8'b1111_1110;
		Dminus[64] = 8'b1111_1111;
		Dminus[65] = 8'b1111_1111;
		Dminus[66] = 8'b1111_1111;
		Dminus[67] = 8'b1111_1111;
		Dminus[68] = 8'b1111_1111;
		Dminus[69] = 8'b1111_1111;
		Dminus[70] = 8'b1111_1111;
		Dminus[71] = 8'b1111_1111;
		Dminus[72] = 8'b1111_1111;
		Dminus[73] = 8'b1111_1111;
		Dminus[74] = 8'b1111_1111;
		Dminus[75] = 8'b1111_1111;
		Dminus[76] = 8'b1111_1111;
		Dminus[77] = 8'b1111_1111;
		Dminus[78] = 8'b1111_1111;
		Dminus[79] = 8'b1111_1111;
		Dminus[80] = 8'b1111_1111;
		Dminus[81] = 8'b1111_1111;
		Dminus[82] = 8'b1111_1111;
		Dminus[83] = 8'b1111_1111;
		Dminus[84] = 8'b1111_1111;
		Dminus[85] = 8'b1111_1111;
		Dminus[86] = 8'b1111_1111;
		Dminus[87] = 8'b1111_1111;
		Dminus[88] = 8'b1111_1111;
		Dminus[89] = 8'b0000_0000;
		Dminus[90] = 8'b0000_0000;
		Dminus[91] = 8'b0000_0000;
		Dminus[92] = 8'b0000_0000;
		Dminus[93] = 8'b0000_0000;
		Dminus[94] = 8'b0000_0000;
		Dminus[95] = 8'b0000_0000;
		Dminus[96] = 8'b0000_0000;
		Dminus[97] = 8'b0000_0000;
		Dminus[98] = 8'b0000_0000;
		Dminus[99] = 8'b0000_0000;
		Dminus[100] = 8'b0000_0000;
		Dminus[101] = 8'b0000_0000;
		Dminus[102] = 8'b0000_0000;
		Dminus[103] = 8'b0000_0000;
		Dminus[104] = 8'b0000_0000;
		Dminus[105] = 8'b0000_0000;
		Dminus[106] = 8'b0000_0000;
		Dminus[107] = 8'b0000_0000;
		Dminus[108] = 8'b0000_0000;
		Dminus[109] = 8'b0000_0000;
		Dminus[110] = 8'b0000_0000;
		Dminus[111] = 8'b0000_0000;
		Dminus[112] = 8'b0000_0000;
		Dminus[113] = 8'b0000_0000;
		Dminus[114] = 8'b0000_0000;
		Dminus[115] = 8'b0000_0000;
		Dminus[116] = 8'b0000_0000;
		Dminus[117] = 8'b0000_0000;
		Dminus[118] = 8'b0000_0000;
		Dminus[119] = 8'b0000_0000;
		Dminus[120] = 8'b0000_0000;
		Dminus[121] = 8'b0000_0000;
		Dminus[122] = 8'b0000_0000;
		Dminus[123] = 8'b0000_0000;
		Dminus[124] = 8'b0000_0000;
		Dminus[125] = 8'b0000_0000;
		Dminus[126] = 8'b0000_0000;
		Dminus[127] = 8'b0000_0000;
		Dplus[1] = 8'b0001_0000;
		Dplus[2] = 8'b0000_1111;
		Dplus[3] = 8'b0000_1111;
		Dplus[4] = 8'b0000_1110;
		Dplus[5] = 8'b0000_1110;
		Dplus[6] = 8'b0000_1101;
		Dplus[7] = 8'b0000_1101;
		Dplus[8] = 8'b0000_1100;
		Dplus[9] = 8'b0000_1100;
		Dplus[10] = 8'b0000_1100;
		Dplus[11] = 8'b0000_1011;
		Dplus[12] = 8'b0000_1011;
		Dplus[13] = 8'b0000_1010;
		Dplus[14] = 8'b0000_1010;
		Dplus[15] = 8'b0000_1010;
		Dplus[16] = 8'b0000_1001;
		Dplus[17] = 8'b0000_1001;
		Dplus[18] = 8'b0000_1001;
		Dplus[19] = 8'b0000_1000;
		Dplus[20] = 8'b0000_1000;
		Dplus[21] = 8'b0000_1000;
		Dplus[22] = 8'b0000_1000;
		Dplus[23] = 8'b0000_0111;
		Dplus[24] = 8'b0000_0111;
		Dplus[25] = 8'b0000_0111;
		Dplus[26] = 8'b0000_0110;
		Dplus[27] = 8'b0000_0110;
		Dplus[28] = 8'b0000_0110;
		Dplus[29] = 8'b0000_0110;
		Dplus[30] = 8'b0000_0110;
		Dplus[31] = 8'b0000_0101;
		Dplus[32] = 8'b0000_0101;
		Dplus[33] = 8'b0000_0101;
		Dplus[34] = 8'b0000_0101;
		Dplus[35] = 8'b0000_0101;
		Dplus[36] = 8'b0000_0100;
		Dplus[37] = 8'b0000_0100;
		Dplus[38] = 8'b0000_0100;
		Dplus[39] = 8'b0000_0100;
		Dplus[40] = 8'b0000_0100;
		Dplus[41] = 8'b0000_0100;
		Dplus[42] = 8'b0000_0011;
		Dplus[43] = 8'b0000_0011;
		Dplus[44] = 8'b0000_0011;
		Dplus[45] = 8'b0000_0011;
		Dplus[46] = 8'b0000_0011;
		Dplus[47] = 8'b0000_0011;
		Dplus[48] = 8'b0000_0011;
		Dplus[49] = 8'b0000_0011;
		Dplus[50] = 8'b0000_0011;
		Dplus[51] = 8'b0000_0010;
		Dplus[52] = 8'b0000_0010;
		Dplus[53] = 8'b0000_0010;
		Dplus[54] = 8'b0000_0010;
		Dplus[55] = 8'b0000_0010;
		Dplus[56] = 8'b0000_0010;
		Dplus[57] = 8'b0000_0010;
		Dplus[58] = 8'b0000_0010;
		Dplus[59] = 8'b0000_0010;
		Dplus[60] = 8'b0000_0010;
		Dplus[61] = 8'b0000_0010;
		Dplus[62] = 8'b0000_0010;
		Dplus[63] = 8'b0000_0001;
		Dplus[64] = 8'b0000_0001;
		Dplus[65] = 8'b0000_0001;
		Dplus[66] = 8'b0000_0001;
		Dplus[67] = 8'b0000_0001;
		Dplus[68] = 8'b0000_0001;
		Dplus[69] = 8'b0000_0001;
		Dplus[70] = 8'b0000_0001;
		Dplus[71] = 8'b0000_0001;
		Dplus[72] = 8'b0000_0001;
		Dplus[73] = 8'b0000_0001;
		Dplus[74] = 8'b0000_0001;
		Dplus[75] = 8'b0000_0001;
		Dplus[76] = 8'b0000_0001;
		Dplus[77] = 8'b0000_0001;
		Dplus[78] = 8'b0000_0001;
		Dplus[79] = 8'b0000_0001;
		Dplus[80] = 8'b0000_0001;
		Dplus[81] = 8'b0000_0001;
		Dplus[82] = 8'b0000_0001;
		Dplus[83] = 8'b0000_0001;
		Dplus[84] = 8'b0000_0001;
		Dplus[85] = 8'b0000_0001;
		Dplus[86] = 8'b0000_0001;
		Dplus[87] = 8'b0000_0001;
		Dplus[88] = 8'b0000_0001;
		Dplus[89] = 8'b0000_0000;
		Dplus[90] = 8'b0000_0000;
		Dplus[91] = 8'b0000_0000;
		Dplus[92] = 8'b0000_0000;
		Dplus[93] = 8'b0000_0000;
		Dplus[94] = 8'b0000_0000;
		Dplus[95] = 8'b0000_0000;
		Dplus[96] = 8'b0000_0000;
		Dplus[97] = 8'b0000_0000;
		Dplus[98] = 8'b0000_0000;
		Dplus[99] = 8'b0000_0000;
		Dplus[100] = 8'b0000_0000;
		Dplus[101] = 8'b0000_0000;
		Dplus[102] = 8'b0000_0000;
		Dplus[103] = 8'b0000_0000;
		Dplus[104] = 8'b0000_0000;
		Dplus[105] = 8'b0000_0000;
		Dplus[106] = 8'b0000_0000;
		Dplus[107] = 8'b0000_0000;
		Dplus[108] = 8'b0000_0000;
		Dplus[109] = 8'b0000_0000;
		Dplus[110] = 8'b0000_0000;
		Dplus[111] = 8'b0000_0000;
		Dplus[112] = 8'b0000_0000;
		Dplus[113] = 8'b0000_0000;
		Dplus[114] = 8'b0000_0000;
		Dplus[115] = 8'b0000_0000;
		Dplus[116] = 8'b0000_0000;
		Dplus[117] = 8'b0000_0000;
		Dplus[118] = 8'b0000_0000;
		Dplus[119] = 8'b0000_0000;
		Dplus[120] = 8'b0000_0000;
		Dplus[121] = 8'b0000_0000;
		Dplus[122] = 8'b0000_0000;
		Dplus[123] = 8'b0000_0000;
		Dplus[124] = 8'b0000_0000;
		Dplus[125] = 8'b0000_0000;
		Dplus[126] = 8'b0000_0000;
		Dplus[127] = 8'b0000_0000;
end
endmodule
