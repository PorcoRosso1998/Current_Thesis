module Tables();
	reg [5:0] Dplus[63:0];
	reg [5:0] Dminus[63:0];
	reg [4:0] DminusInteger[15:0];
	reg [4:0] DplusInteger[15:0];
	initial begin
		Dminus[1] = 10'b11010_01111;
		Dminus[2] = 10'b11011_01110;
		Dminus[3] = 10'b11100_00000;
		Dminus[4] = 10'b11100_01101;
		Dminus[5] = 10'b11100_10111;
		Dminus[6] = 10'b11100_11111;
		Dminus[7] = 10'b11101_00101;
		Dminus[8] = 10'b11101_01011;
		Dminus[9] = 10'b11101_10000;
		Dminus[10] = 10'b11101_10100;
		Dminus[11] = 10'b11101_11000;
		Dminus[12] = 10'b11101_11100;
		Dminus[13] = 10'b11101_11111;
		Dminus[14] = 10'b11110_00010;
		Dminus[15] = 10'b11110_00101;
		Dminus[16] = 10'b11110_00111;
		Dminus[17] = 10'b11110_01010;
		Dminus[18] = 10'b11110_01100;
		Dminus[19] = 10'b11110_01110;
		Dminus[20] = 10'b11110_10000;
		Dminus[21] = 10'b11110_10010;
		Dminus[22] = 10'b11110_10011;
		Dminus[23] = 10'b11110_10101;
		Dminus[24] = 10'b11110_10110;
		Dminus[25] = 10'b11110_11000;
		Dminus[26] = 10'b11110_11001;
		Dminus[27] = 10'b11110_11010;
		Dminus[28] = 10'b11110_11100;
		Dminus[29] = 10'b11110_11101;
		Dminus[30] = 10'b11110_11110;
		Dminus[31] = 10'b11110_11111;
		Dminus[32] = 10'b11111_00000;
		Dminus[33] = 10'b11111_00001;
		Dminus[34] = 10'b11111_00010;
		Dminus[35] = 10'b11111_00011;
		Dminus[36] = 10'b11111_00100;
		Dminus[37] = 10'b11111_00101;
		Dminus[38] = 10'b11111_00101;
		Dminus[39] = 10'b11111_00110;
		Dminus[40] = 10'b11111_00111;
		Dminus[41] = 10'b11111_01000;
		Dminus[42] = 10'b11111_01000;
		Dminus[43] = 10'b11111_01001;
		Dminus[44] = 10'b11111_01010;
		Dminus[45] = 10'b11111_01010;
		Dminus[46] = 10'b11111_01011;
		Dminus[47] = 10'b11111_01011;
		Dminus[48] = 10'b11111_01100;
		Dminus[49] = 10'b11111_01100;
		Dminus[50] = 10'b11111_01101;
		Dminus[51] = 10'b11111_01101;
		Dminus[52] = 10'b11111_01110;
		Dminus[53] = 10'b11111_01110;
		Dminus[54] = 10'b11111_01111;
		Dminus[55] = 10'b11111_01111;
		Dminus[56] = 10'b11111_10000;
		Dminus[57] = 10'b11111_10000;
		Dminus[58] = 10'b11111_10001;
		Dminus[59] = 10'b11111_10001;
		Dminus[60] = 10'b11111_10001;
		Dminus[61] = 10'b11111_10010;
		Dminus[62] = 10'b11111_10010;
		Dminus[63] = 10'b11111_10010;
		Dplus[1] = 10'b00001_00000;
		Dplus[2] = 10'b00000_11111;
		Dplus[3] = 10'b00000_11111;
		Dplus[4] = 10'b00000_11110;
		Dplus[5] = 10'b00000_11110;
		Dplus[6] = 10'b00000_11101;
		Dplus[7] = 10'b00000_11101;
		Dplus[8] = 10'b00000_11100;
		Dplus[9] = 10'b00000_11100;
		Dplus[10] = 10'b00000_11011;
		Dplus[11] = 10'b00000_11011;
		Dplus[12] = 10'b00000_11010;
		Dplus[13] = 10'b00000_11010;
		Dplus[14] = 10'b00000_11010;
		Dplus[15] = 10'b00000_11001;
		Dplus[16] = 10'b00000_11001;
		Dplus[17] = 10'b00000_11000;
		Dplus[18] = 10'b00000_11000;
		Dplus[19] = 10'b00000_10111;
		Dplus[20] = 10'b00000_10111;
		Dplus[21] = 10'b00000_10111;
		Dplus[22] = 10'b00000_10110;
		Dplus[23] = 10'b00000_10110;
		Dplus[24] = 10'b00000_10110;
		Dplus[25] = 10'b00000_10101;
		Dplus[26] = 10'b00000_10101;
		Dplus[27] = 10'b00000_10100;
		Dplus[28] = 10'b00000_10100;
		Dplus[29] = 10'b00000_10100;
		Dplus[30] = 10'b00000_10011;
		Dplus[31] = 10'b00000_10011;
		Dplus[32] = 10'b00000_10011;
		Dplus[33] = 10'b00000_10010;
		Dplus[34] = 10'b00000_10010;
		Dplus[35] = 10'b00000_10010;
		Dplus[36] = 10'b00000_10001;
		Dplus[37] = 10'b00000_10001;
		Dplus[38] = 10'b00000_10001;
		Dplus[39] = 10'b00000_10001;
		Dplus[40] = 10'b00000_10000;
		Dplus[41] = 10'b00000_10000;
		Dplus[42] = 10'b00000_10000;
		Dplus[43] = 10'b00000_01111;
		Dplus[44] = 10'b00000_01111;
		Dplus[45] = 10'b00000_01111;
		Dplus[46] = 10'b00000_01111;
		Dplus[47] = 10'b00000_01110;
		Dplus[48] = 10'b00000_01110;
		Dplus[49] = 10'b00000_01110;
		Dplus[50] = 10'b00000_01101;
		Dplus[51] = 10'b00000_01101;
		Dplus[52] = 10'b00000_01101;
		Dplus[53] = 10'b00000_01101;
		Dplus[54] = 10'b00000_01100;
		Dplus[55] = 10'b00000_01100;
		Dplus[56] = 10'b00000_01100;
		Dplus[57] = 10'b00000_01100;
		Dplus[58] = 10'b00000_01100;
		Dplus[59] = 10'b00000_01011;
		Dplus[60] = 10'b00000_01011;
		Dplus[61] = 10'b00000_01011;
		Dplus[62] = 10'b00000_01011;
		Dplus[63] = 10'b00000_01011;
		Dplus[2] = 10'b00000_01010;
		Dplus[3] = 10'b00000_00101;
		Dplus[4] = 10'b00000_00011;
		Dplus[5] = 10'b00000_00001;
		Dplus[6] = 10'b00000_00001;
		Dplus[7] = 10'b00000_00000;
		Dplus[8] = 10'b00000_00000;
		Dplus[9] = 10'b00000_00000;
		Dplus[10] = 10'b00000_00000;
		Dplus[11] = 10'b00000_00000;
		Dplus[12] = 10'b00000_00000;
		Dplus[13] = 10'b00000_00000;
		Dplus[14] = 10'b00000_00000;
		Dplus[15] = 10'b00000_00000;
		Dminus[2] = 10'b11111_10011;
		Dminus[3] = 10'b11111_11010;
		Dminus[4] = 10'b11111_11101;
		Dminus[5] = 10'b11111_11111;
		Dminus[6] = 10'b11111_11111;
		Dminus[7] = 10'b00000_00000;
		Dminus[8] = 10'b00000_00000;
		Dminus[9] = 10'b00000_00000;
		Dminus[10] = 10'b00000_00000;
		Dminus[11] = 10'b00000_00000;
		Dminus[12] = 10'b00000_00000;
		Dminus[13] = 10'b00000_00000;
		Dminus[14] = 10'b00000_00000;
		Dminus[15] = 10'b00000_00000;
end
endmodule
