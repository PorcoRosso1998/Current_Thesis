module Tables();
	reg [11:0] logarithm_table[2047:0];
	reg [11:0] Dplus[2047:0];
	reg [11:0] Dminus[2047:0];
	initial begin
		logarithm_table[1] = 12'b111010_000000;
		logarithm_table[2] = 12'b111011_000000;
		logarithm_table[3] = 12'b111011_100101;
		logarithm_table[4] = 12'b111100_000000;
		logarithm_table[5] = 12'b111100_010101;
		logarithm_table[6] = 12'b111100_100101;
		logarithm_table[7] = 12'b111100_110100;
		logarithm_table[8] = 12'b111101_000000;
		logarithm_table[9] = 12'b111101_001011;
		logarithm_table[10] = 12'b111101_010101;
		logarithm_table[11] = 12'b111101_011101;
		logarithm_table[12] = 12'b111101_100101;
		logarithm_table[13] = 12'b111101_101101;
		logarithm_table[14] = 12'b111101_110100;
		logarithm_table[15] = 12'b111101_111010;
		logarithm_table[16] = 12'b111110_000000;
		logarithm_table[17] = 12'b111110_000110;
		logarithm_table[18] = 12'b111110_001011;
		logarithm_table[19] = 12'b111110_010000;
		logarithm_table[20] = 12'b111110_010101;
		logarithm_table[21] = 12'b111110_011001;
		logarithm_table[22] = 12'b111110_011101;
		logarithm_table[23] = 12'b111110_100010;
		logarithm_table[24] = 12'b111110_100101;
		logarithm_table[25] = 12'b111110_101001;
		logarithm_table[26] = 12'b111110_101101;
		logarithm_table[27] = 12'b111110_110000;
		logarithm_table[28] = 12'b111110_110100;
		logarithm_table[29] = 12'b111110_110111;
		logarithm_table[30] = 12'b111110_111010;
		logarithm_table[31] = 12'b111110_111101;
		logarithm_table[32] = 12'b111111_000000;
		logarithm_table[33] = 12'b111111_000011;
		logarithm_table[34] = 12'b111111_000110;
		logarithm_table[35] = 12'b111111_001000;
		logarithm_table[36] = 12'b111111_001011;
		logarithm_table[37] = 12'b111111_001101;
		logarithm_table[38] = 12'b111111_010000;
		logarithm_table[39] = 12'b111111_010010;
		logarithm_table[40] = 12'b111111_010101;
		logarithm_table[41] = 12'b111111_010111;
		logarithm_table[42] = 12'b111111_011001;
		logarithm_table[43] = 12'b111111_011011;
		logarithm_table[44] = 12'b111111_011101;
		logarithm_table[45] = 12'b111111_011111;
		logarithm_table[46] = 12'b111111_100010;
		logarithm_table[47] = 12'b111111_100011;
		logarithm_table[48] = 12'b111111_100101;
		logarithm_table[49] = 12'b111111_100111;
		logarithm_table[50] = 12'b111111_101001;
		logarithm_table[51] = 12'b111111_101011;
		logarithm_table[52] = 12'b111111_101101;
		logarithm_table[53] = 12'b111111_101111;
		logarithm_table[54] = 12'b111111_110000;
		logarithm_table[55] = 12'b111111_110010;
		logarithm_table[56] = 12'b111111_110100;
		logarithm_table[57] = 12'b111111_110101;
		logarithm_table[58] = 12'b111111_110111;
		logarithm_table[59] = 12'b111111_111000;
		logarithm_table[60] = 12'b111111_111010;
		logarithm_table[61] = 12'b111111_111100;
		logarithm_table[62] = 12'b111111_111101;
		logarithm_table[63] = 12'b111111_111111;
		logarithm_table[64] = 12'b000000_000000;
		logarithm_table[65] = 12'b000000_000001;
		logarithm_table[66] = 12'b000000_000011;
		logarithm_table[67] = 12'b000000_000100;
		logarithm_table[68] = 12'b000000_000110;
		logarithm_table[69] = 12'b000000_000111;
		logarithm_table[70] = 12'b000000_001000;
		logarithm_table[71] = 12'b000000_001010;
		logarithm_table[72] = 12'b000000_001011;
		logarithm_table[73] = 12'b000000_001100;
		logarithm_table[74] = 12'b000000_001101;
		logarithm_table[75] = 12'b000000_001111;
		logarithm_table[76] = 12'b000000_010000;
		logarithm_table[77] = 12'b000000_010001;
		logarithm_table[78] = 12'b000000_010010;
		logarithm_table[79] = 12'b000000_010011;
		logarithm_table[80] = 12'b000000_010101;
		logarithm_table[81] = 12'b000000_010110;
		logarithm_table[82] = 12'b000000_010111;
		logarithm_table[83] = 12'b000000_011000;
		logarithm_table[84] = 12'b000000_011001;
		logarithm_table[85] = 12'b000000_011010;
		logarithm_table[86] = 12'b000000_011011;
		logarithm_table[87] = 12'b000000_011100;
		logarithm_table[88] = 12'b000000_011101;
		logarithm_table[89] = 12'b000000_011110;
		logarithm_table[90] = 12'b000000_011111;
		logarithm_table[91] = 12'b000000_100000;
		logarithm_table[92] = 12'b000000_100010;
		logarithm_table[93] = 12'b000000_100011;
		logarithm_table[94] = 12'b000000_100011;
		logarithm_table[95] = 12'b000000_100100;
		logarithm_table[96] = 12'b000000_100101;
		logarithm_table[97] = 12'b000000_100110;
		logarithm_table[98] = 12'b000000_100111;
		logarithm_table[99] = 12'b000000_101000;
		logarithm_table[100] = 12'b000000_101001;
		logarithm_table[101] = 12'b000000_101010;
		logarithm_table[102] = 12'b000000_101011;
		logarithm_table[103] = 12'b000000_101100;
		logarithm_table[104] = 12'b000000_101101;
		logarithm_table[105] = 12'b000000_101110;
		logarithm_table[106] = 12'b000000_101111;
		logarithm_table[107] = 12'b000000_101111;
		logarithm_table[108] = 12'b000000_110000;
		logarithm_table[109] = 12'b000000_110001;
		logarithm_table[110] = 12'b000000_110010;
		logarithm_table[111] = 12'b000000_110011;
		logarithm_table[112] = 12'b000000_110100;
		logarithm_table[113] = 12'b000000_110100;
		logarithm_table[114] = 12'b000000_110101;
		logarithm_table[115] = 12'b000000_110110;
		logarithm_table[116] = 12'b000000_110111;
		logarithm_table[117] = 12'b000000_111000;
		logarithm_table[118] = 12'b000000_111000;
		logarithm_table[119] = 12'b000000_111001;
		logarithm_table[120] = 12'b000000_111010;
		logarithm_table[121] = 12'b000000_111011;
		logarithm_table[122] = 12'b000000_111100;
		logarithm_table[123] = 12'b000000_111100;
		logarithm_table[124] = 12'b000000_111101;
		logarithm_table[125] = 12'b000000_111110;
		logarithm_table[126] = 12'b000000_111111;
		logarithm_table[127] = 12'b000000_111111;
		logarithm_table[128] = 12'b000001_000000;
		logarithm_table[129] = 12'b000001_000001;
		logarithm_table[130] = 12'b000001_000001;
		logarithm_table[131] = 12'b000001_000010;
		logarithm_table[132] = 12'b000001_000011;
		logarithm_table[133] = 12'b000001_000100;
		logarithm_table[134] = 12'b000001_000100;
		logarithm_table[135] = 12'b000001_000101;
		logarithm_table[136] = 12'b000001_000110;
		logarithm_table[137] = 12'b000001_000110;
		logarithm_table[138] = 12'b000001_000111;
		logarithm_table[139] = 12'b000001_001000;
		logarithm_table[140] = 12'b000001_001000;
		logarithm_table[141] = 12'b000001_001001;
		logarithm_table[142] = 12'b000001_001010;
		logarithm_table[143] = 12'b000001_001010;
		logarithm_table[144] = 12'b000001_001011;
		logarithm_table[145] = 12'b000001_001100;
		logarithm_table[146] = 12'b000001_001100;
		logarithm_table[147] = 12'b000001_001101;
		logarithm_table[148] = 12'b000001_001101;
		logarithm_table[149] = 12'b000001_001110;
		logarithm_table[150] = 12'b000001_001111;
		logarithm_table[151] = 12'b000001_001111;
		logarithm_table[152] = 12'b000001_010000;
		logarithm_table[153] = 12'b000001_010000;
		logarithm_table[154] = 12'b000001_010001;
		logarithm_table[155] = 12'b000001_010010;
		logarithm_table[156] = 12'b000001_010010;
		logarithm_table[157] = 12'b000001_010011;
		logarithm_table[158] = 12'b000001_010011;
		logarithm_table[159] = 12'b000001_010100;
		logarithm_table[160] = 12'b000001_010101;
		logarithm_table[161] = 12'b000001_010101;
		logarithm_table[162] = 12'b000001_010110;
		logarithm_table[163] = 12'b000001_010110;
		logarithm_table[164] = 12'b000001_010111;
		logarithm_table[165] = 12'b000001_010111;
		logarithm_table[166] = 12'b000001_011000;
		logarithm_table[167] = 12'b000001_011001;
		logarithm_table[168] = 12'b000001_011001;
		logarithm_table[169] = 12'b000001_011010;
		logarithm_table[170] = 12'b000001_011010;
		logarithm_table[171] = 12'b000001_011011;
		logarithm_table[172] = 12'b000001_011011;
		logarithm_table[173] = 12'b000001_011100;
		logarithm_table[174] = 12'b000001_011100;
		logarithm_table[175] = 12'b000001_011101;
		logarithm_table[176] = 12'b000001_011101;
		logarithm_table[177] = 12'b000001_011110;
		logarithm_table[178] = 12'b000001_011110;
		logarithm_table[179] = 12'b000001_011111;
		logarithm_table[180] = 12'b000001_011111;
		logarithm_table[181] = 12'b000001_100000;
		logarithm_table[182] = 12'b000001_100000;
		logarithm_table[183] = 12'b000001_100001;
		logarithm_table[184] = 12'b000001_100010;
		logarithm_table[185] = 12'b000001_100010;
		logarithm_table[186] = 12'b000001_100011;
		logarithm_table[187] = 12'b000001_100011;
		logarithm_table[188] = 12'b000001_100011;
		logarithm_table[189] = 12'b000001_100100;
		logarithm_table[190] = 12'b000001_100100;
		logarithm_table[191] = 12'b000001_100101;
		logarithm_table[192] = 12'b000001_100101;
		logarithm_table[193] = 12'b000001_100110;
		logarithm_table[194] = 12'b000001_100110;
		logarithm_table[195] = 12'b000001_100111;
		logarithm_table[196] = 12'b000001_100111;
		logarithm_table[197] = 12'b000001_101000;
		logarithm_table[198] = 12'b000001_101000;
		logarithm_table[199] = 12'b000001_101001;
		logarithm_table[200] = 12'b000001_101001;
		logarithm_table[201] = 12'b000001_101010;
		logarithm_table[202] = 12'b000001_101010;
		logarithm_table[203] = 12'b000001_101011;
		logarithm_table[204] = 12'b000001_101011;
		logarithm_table[205] = 12'b000001_101011;
		logarithm_table[206] = 12'b000001_101100;
		logarithm_table[207] = 12'b000001_101100;
		logarithm_table[208] = 12'b000001_101101;
		logarithm_table[209] = 12'b000001_101101;
		logarithm_table[210] = 12'b000001_101110;
		logarithm_table[211] = 12'b000001_101110;
		logarithm_table[212] = 12'b000001_101111;
		logarithm_table[213] = 12'b000001_101111;
		logarithm_table[214] = 12'b000001_101111;
		logarithm_table[215] = 12'b000001_110000;
		logarithm_table[216] = 12'b000001_110000;
		logarithm_table[217] = 12'b000001_110001;
		logarithm_table[218] = 12'b000001_110001;
		logarithm_table[219] = 12'b000001_110010;
		logarithm_table[220] = 12'b000001_110010;
		logarithm_table[221] = 12'b000001_110010;
		logarithm_table[222] = 12'b000001_110011;
		logarithm_table[223] = 12'b000001_110011;
		logarithm_table[224] = 12'b000001_110100;
		logarithm_table[225] = 12'b000001_110100;
		logarithm_table[226] = 12'b000001_110100;
		logarithm_table[227] = 12'b000001_110101;
		logarithm_table[228] = 12'b000001_110101;
		logarithm_table[229] = 12'b000001_110110;
		logarithm_table[230] = 12'b000001_110110;
		logarithm_table[231] = 12'b000001_110111;
		logarithm_table[232] = 12'b000001_110111;
		logarithm_table[233] = 12'b000001_110111;
		logarithm_table[234] = 12'b000001_111000;
		logarithm_table[235] = 12'b000001_111000;
		logarithm_table[236] = 12'b000001_111000;
		logarithm_table[237] = 12'b000001_111001;
		logarithm_table[238] = 12'b000001_111001;
		logarithm_table[239] = 12'b000001_111010;
		logarithm_table[240] = 12'b000001_111010;
		logarithm_table[241] = 12'b000001_111010;
		logarithm_table[242] = 12'b000001_111011;
		logarithm_table[243] = 12'b000001_111011;
		logarithm_table[244] = 12'b000001_111100;
		logarithm_table[245] = 12'b000001_111100;
		logarithm_table[246] = 12'b000001_111100;
		logarithm_table[247] = 12'b000001_111101;
		logarithm_table[248] = 12'b000001_111101;
		logarithm_table[249] = 12'b000001_111101;
		logarithm_table[250] = 12'b000001_111110;
		logarithm_table[251] = 12'b000001_111110;
		logarithm_table[252] = 12'b000001_111111;
		logarithm_table[253] = 12'b000001_111111;
		logarithm_table[254] = 12'b000001_111111;
		logarithm_table[255] = 12'b000010_000000;
		logarithm_table[256] = 12'b000010_000000;
		logarithm_table[257] = 12'b000010_000000;
		logarithm_table[258] = 12'b000010_000001;
		logarithm_table[259] = 12'b000010_000001;
		logarithm_table[260] = 12'b000010_000001;
		logarithm_table[261] = 12'b000010_000010;
		logarithm_table[262] = 12'b000010_000010;
		logarithm_table[263] = 12'b000010_000010;
		logarithm_table[264] = 12'b000010_000011;
		logarithm_table[265] = 12'b000010_000011;
		logarithm_table[266] = 12'b000010_000100;
		logarithm_table[267] = 12'b000010_000100;
		logarithm_table[268] = 12'b000010_000100;
		logarithm_table[269] = 12'b000010_000101;
		logarithm_table[270] = 12'b000010_000101;
		logarithm_table[271] = 12'b000010_000101;
		logarithm_table[272] = 12'b000010_000110;
		logarithm_table[273] = 12'b000010_000110;
		logarithm_table[274] = 12'b000010_000110;
		logarithm_table[275] = 12'b000010_000111;
		logarithm_table[276] = 12'b000010_000111;
		logarithm_table[277] = 12'b000010_000111;
		logarithm_table[278] = 12'b000010_001000;
		logarithm_table[279] = 12'b000010_001000;
		logarithm_table[280] = 12'b000010_001000;
		logarithm_table[281] = 12'b000010_001001;
		logarithm_table[282] = 12'b000010_001001;
		logarithm_table[283] = 12'b000010_001001;
		logarithm_table[284] = 12'b000010_001010;
		logarithm_table[285] = 12'b000010_001010;
		logarithm_table[286] = 12'b000010_001010;
		logarithm_table[287] = 12'b000010_001011;
		logarithm_table[288] = 12'b000010_001011;
		logarithm_table[289] = 12'b000010_001011;
		logarithm_table[290] = 12'b000010_001100;
		logarithm_table[291] = 12'b000010_001100;
		logarithm_table[292] = 12'b000010_001100;
		logarithm_table[293] = 12'b000010_001100;
		logarithm_table[294] = 12'b000010_001101;
		logarithm_table[295] = 12'b000010_001101;
		logarithm_table[296] = 12'b000010_001101;
		logarithm_table[297] = 12'b000010_001110;
		logarithm_table[298] = 12'b000010_001110;
		logarithm_table[299] = 12'b000010_001110;
		logarithm_table[300] = 12'b000010_001111;
		logarithm_table[301] = 12'b000010_001111;
		logarithm_table[302] = 12'b000010_001111;
		logarithm_table[303] = 12'b000010_010000;
		logarithm_table[304] = 12'b000010_010000;
		logarithm_table[305] = 12'b000010_010000;
		logarithm_table[306] = 12'b000010_010000;
		logarithm_table[307] = 12'b000010_010001;
		logarithm_table[308] = 12'b000010_010001;
		logarithm_table[309] = 12'b000010_010001;
		logarithm_table[310] = 12'b000010_010010;
		logarithm_table[311] = 12'b000010_010010;
		logarithm_table[312] = 12'b000010_010010;
		logarithm_table[313] = 12'b000010_010011;
		logarithm_table[314] = 12'b000010_010011;
		logarithm_table[315] = 12'b000010_010011;
		logarithm_table[316] = 12'b000010_010011;
		logarithm_table[317] = 12'b000010_010100;
		logarithm_table[318] = 12'b000010_010100;
		logarithm_table[319] = 12'b000010_010100;
		logarithm_table[320] = 12'b000010_010101;
		logarithm_table[321] = 12'b000010_010101;
		logarithm_table[322] = 12'b000010_010101;
		logarithm_table[323] = 12'b000010_010101;
		logarithm_table[324] = 12'b000010_010110;
		logarithm_table[325] = 12'b000010_010110;
		logarithm_table[326] = 12'b000010_010110;
		logarithm_table[327] = 12'b000010_010111;
		logarithm_table[328] = 12'b000010_010111;
		logarithm_table[329] = 12'b000010_010111;
		logarithm_table[330] = 12'b000010_010111;
		logarithm_table[331] = 12'b000010_011000;
		logarithm_table[332] = 12'b000010_011000;
		logarithm_table[333] = 12'b000010_011000;
		logarithm_table[334] = 12'b000010_011001;
		logarithm_table[335] = 12'b000010_011001;
		logarithm_table[336] = 12'b000010_011001;
		logarithm_table[337] = 12'b000010_011001;
		logarithm_table[338] = 12'b000010_011010;
		logarithm_table[339] = 12'b000010_011010;
		logarithm_table[340] = 12'b000010_011010;
		logarithm_table[341] = 12'b000010_011010;
		logarithm_table[342] = 12'b000010_011011;
		logarithm_table[343] = 12'b000010_011011;
		logarithm_table[344] = 12'b000010_011011;
		logarithm_table[345] = 12'b000010_011100;
		logarithm_table[346] = 12'b000010_011100;
		logarithm_table[347] = 12'b000010_011100;
		logarithm_table[348] = 12'b000010_011100;
		logarithm_table[349] = 12'b000010_011101;
		logarithm_table[350] = 12'b000010_011101;
		logarithm_table[351] = 12'b000010_011101;
		logarithm_table[352] = 12'b000010_011101;
		logarithm_table[353] = 12'b000010_011110;
		logarithm_table[354] = 12'b000010_011110;
		logarithm_table[355] = 12'b000010_011110;
		logarithm_table[356] = 12'b000010_011110;
		logarithm_table[357] = 12'b000010_011111;
		logarithm_table[358] = 12'b000010_011111;
		logarithm_table[359] = 12'b000010_011111;
		logarithm_table[360] = 12'b000010_011111;
		logarithm_table[361] = 12'b000010_100000;
		logarithm_table[362] = 12'b000010_100000;
		logarithm_table[363] = 12'b000010_100000;
		logarithm_table[364] = 12'b000010_100000;
		logarithm_table[365] = 12'b000010_100001;
		logarithm_table[366] = 12'b000010_100001;
		logarithm_table[367] = 12'b000010_100001;
		logarithm_table[368] = 12'b000010_100010;
		logarithm_table[369] = 12'b000010_100010;
		logarithm_table[370] = 12'b000010_100010;
		logarithm_table[371] = 12'b000010_100010;
		logarithm_table[372] = 12'b000010_100011;
		logarithm_table[373] = 12'b000010_100011;
		logarithm_table[374] = 12'b000010_100011;
		logarithm_table[375] = 12'b000010_100011;
		logarithm_table[376] = 12'b000010_100011;
		logarithm_table[377] = 12'b000010_100100;
		logarithm_table[378] = 12'b000010_100100;
		logarithm_table[379] = 12'b000010_100100;
		logarithm_table[380] = 12'b000010_100100;
		logarithm_table[381] = 12'b000010_100101;
		logarithm_table[382] = 12'b000010_100101;
		logarithm_table[383] = 12'b000010_100101;
		logarithm_table[384] = 12'b000010_100101;
		logarithm_table[385] = 12'b000010_100110;
		logarithm_table[386] = 12'b000010_100110;
		logarithm_table[387] = 12'b000010_100110;
		logarithm_table[388] = 12'b000010_100110;
		logarithm_table[389] = 12'b000010_100111;
		logarithm_table[390] = 12'b000010_100111;
		logarithm_table[391] = 12'b000010_100111;
		logarithm_table[392] = 12'b000010_100111;
		logarithm_table[393] = 12'b000010_101000;
		logarithm_table[394] = 12'b000010_101000;
		logarithm_table[395] = 12'b000010_101000;
		logarithm_table[396] = 12'b000010_101000;
		logarithm_table[397] = 12'b000010_101001;
		logarithm_table[398] = 12'b000010_101001;
		logarithm_table[399] = 12'b000010_101001;
		logarithm_table[400] = 12'b000010_101001;
		logarithm_table[401] = 12'b000010_101001;
		logarithm_table[402] = 12'b000010_101010;
		logarithm_table[403] = 12'b000010_101010;
		logarithm_table[404] = 12'b000010_101010;
		logarithm_table[405] = 12'b000010_101010;
		logarithm_table[406] = 12'b000010_101011;
		logarithm_table[407] = 12'b000010_101011;
		logarithm_table[408] = 12'b000010_101011;
		logarithm_table[409] = 12'b000010_101011;
		logarithm_table[410] = 12'b000010_101011;
		logarithm_table[411] = 12'b000010_101100;
		logarithm_table[412] = 12'b000010_101100;
		logarithm_table[413] = 12'b000010_101100;
		logarithm_table[414] = 12'b000010_101100;
		logarithm_table[415] = 12'b000010_101101;
		logarithm_table[416] = 12'b000010_101101;
		logarithm_table[417] = 12'b000010_101101;
		logarithm_table[418] = 12'b000010_101101;
		logarithm_table[419] = 12'b000010_101101;
		logarithm_table[420] = 12'b000010_101110;
		logarithm_table[421] = 12'b000010_101110;
		logarithm_table[422] = 12'b000010_101110;
		logarithm_table[423] = 12'b000010_101110;
		logarithm_table[424] = 12'b000010_101111;
		logarithm_table[425] = 12'b000010_101111;
		logarithm_table[426] = 12'b000010_101111;
		logarithm_table[427] = 12'b000010_101111;
		logarithm_table[428] = 12'b000010_101111;
		logarithm_table[429] = 12'b000010_110000;
		logarithm_table[430] = 12'b000010_110000;
		logarithm_table[431] = 12'b000010_110000;
		logarithm_table[432] = 12'b000010_110000;
		logarithm_table[433] = 12'b000010_110001;
		logarithm_table[434] = 12'b000010_110001;
		logarithm_table[435] = 12'b000010_110001;
		logarithm_table[436] = 12'b000010_110001;
		logarithm_table[437] = 12'b000010_110001;
		logarithm_table[438] = 12'b000010_110010;
		logarithm_table[439] = 12'b000010_110010;
		logarithm_table[440] = 12'b000010_110010;
		logarithm_table[441] = 12'b000010_110010;
		logarithm_table[442] = 12'b000010_110010;
		logarithm_table[443] = 12'b000010_110011;
		logarithm_table[444] = 12'b000010_110011;
		logarithm_table[445] = 12'b000010_110011;
		logarithm_table[446] = 12'b000010_110011;
		logarithm_table[447] = 12'b000010_110011;
		logarithm_table[448] = 12'b000010_110100;
		logarithm_table[449] = 12'b000010_110100;
		logarithm_table[450] = 12'b000010_110100;
		logarithm_table[451] = 12'b000010_110100;
		logarithm_table[452] = 12'b000010_110100;
		logarithm_table[453] = 12'b000010_110101;
		logarithm_table[454] = 12'b000010_110101;
		logarithm_table[455] = 12'b000010_110101;
		logarithm_table[456] = 12'b000010_110101;
		logarithm_table[457] = 12'b000010_110110;
		logarithm_table[458] = 12'b000010_110110;
		logarithm_table[459] = 12'b000010_110110;
		logarithm_table[460] = 12'b000010_110110;
		logarithm_table[461] = 12'b000010_110110;
		logarithm_table[462] = 12'b000010_110111;
		logarithm_table[463] = 12'b000010_110111;
		logarithm_table[464] = 12'b000010_110111;
		logarithm_table[465] = 12'b000010_110111;
		logarithm_table[466] = 12'b000010_110111;
		logarithm_table[467] = 12'b000010_111000;
		logarithm_table[468] = 12'b000010_111000;
		logarithm_table[469] = 12'b000010_111000;
		logarithm_table[470] = 12'b000010_111000;
		logarithm_table[471] = 12'b000010_111000;
		logarithm_table[472] = 12'b000010_111000;
		logarithm_table[473] = 12'b000010_111001;
		logarithm_table[474] = 12'b000010_111001;
		logarithm_table[475] = 12'b000010_111001;
		logarithm_table[476] = 12'b000010_111001;
		logarithm_table[477] = 12'b000010_111001;
		logarithm_table[478] = 12'b000010_111010;
		logarithm_table[479] = 12'b000010_111010;
		logarithm_table[480] = 12'b000010_111010;
		logarithm_table[481] = 12'b000010_111010;
		logarithm_table[482] = 12'b000010_111010;
		logarithm_table[483] = 12'b000010_111011;
		logarithm_table[484] = 12'b000010_111011;
		logarithm_table[485] = 12'b000010_111011;
		logarithm_table[486] = 12'b000010_111011;
		logarithm_table[487] = 12'b000010_111011;
		logarithm_table[488] = 12'b000010_111100;
		logarithm_table[489] = 12'b000010_111100;
		logarithm_table[490] = 12'b000010_111100;
		logarithm_table[491] = 12'b000010_111100;
		logarithm_table[492] = 12'b000010_111100;
		logarithm_table[493] = 12'b000010_111101;
		logarithm_table[494] = 12'b000010_111101;
		logarithm_table[495] = 12'b000010_111101;
		logarithm_table[496] = 12'b000010_111101;
		logarithm_table[497] = 12'b000010_111101;
		logarithm_table[498] = 12'b000010_111101;
		logarithm_table[499] = 12'b000010_111110;
		logarithm_table[500] = 12'b000010_111110;
		logarithm_table[501] = 12'b000010_111110;
		logarithm_table[502] = 12'b000010_111110;
		logarithm_table[503] = 12'b000010_111110;
		logarithm_table[504] = 12'b000010_111111;
		logarithm_table[505] = 12'b000010_111111;
		logarithm_table[506] = 12'b000010_111111;
		logarithm_table[507] = 12'b000010_111111;
		logarithm_table[508] = 12'b000010_111111;
		logarithm_table[509] = 12'b000010_111111;
		logarithm_table[510] = 12'b000011_000000;
		logarithm_table[511] = 12'b000011_000000;
		logarithm_table[512] = 12'b000011_000000;
		logarithm_table[513] = 12'b000011_000000;
		logarithm_table[514] = 12'b000011_000000;
		logarithm_table[515] = 12'b000011_000001;
		logarithm_table[516] = 12'b000011_000001;
		logarithm_table[517] = 12'b000011_000001;
		logarithm_table[518] = 12'b000011_000001;
		logarithm_table[519] = 12'b000011_000001;
		logarithm_table[520] = 12'b000011_000001;
		logarithm_table[521] = 12'b000011_000010;
		logarithm_table[522] = 12'b000011_000010;
		logarithm_table[523] = 12'b000011_000010;
		logarithm_table[524] = 12'b000011_000010;
		logarithm_table[525] = 12'b000011_000010;
		logarithm_table[526] = 12'b000011_000010;
		logarithm_table[527] = 12'b000011_000011;
		logarithm_table[528] = 12'b000011_000011;
		logarithm_table[529] = 12'b000011_000011;
		logarithm_table[530] = 12'b000011_000011;
		logarithm_table[531] = 12'b000011_000011;
		logarithm_table[532] = 12'b000011_000100;
		logarithm_table[533] = 12'b000011_000100;
		logarithm_table[534] = 12'b000011_000100;
		logarithm_table[535] = 12'b000011_000100;
		logarithm_table[536] = 12'b000011_000100;
		logarithm_table[537] = 12'b000011_000100;
		logarithm_table[538] = 12'b000011_000101;
		logarithm_table[539] = 12'b000011_000101;
		logarithm_table[540] = 12'b000011_000101;
		logarithm_table[541] = 12'b000011_000101;
		logarithm_table[542] = 12'b000011_000101;
		logarithm_table[543] = 12'b000011_000101;
		logarithm_table[544] = 12'b000011_000110;
		logarithm_table[545] = 12'b000011_000110;
		logarithm_table[546] = 12'b000011_000110;
		logarithm_table[547] = 12'b000011_000110;
		logarithm_table[548] = 12'b000011_000110;
		logarithm_table[549] = 12'b000011_000110;
		logarithm_table[550] = 12'b000011_000111;
		logarithm_table[551] = 12'b000011_000111;
		logarithm_table[552] = 12'b000011_000111;
		logarithm_table[553] = 12'b000011_000111;
		logarithm_table[554] = 12'b000011_000111;
		logarithm_table[555] = 12'b000011_000111;
		logarithm_table[556] = 12'b000011_001000;
		logarithm_table[557] = 12'b000011_001000;
		logarithm_table[558] = 12'b000011_001000;
		logarithm_table[559] = 12'b000011_001000;
		logarithm_table[560] = 12'b000011_001000;
		logarithm_table[561] = 12'b000011_001000;
		logarithm_table[562] = 12'b000011_001001;
		logarithm_table[563] = 12'b000011_001001;
		logarithm_table[564] = 12'b000011_001001;
		logarithm_table[565] = 12'b000011_001001;
		logarithm_table[566] = 12'b000011_001001;
		logarithm_table[567] = 12'b000011_001001;
		logarithm_table[568] = 12'b000011_001010;
		logarithm_table[569] = 12'b000011_001010;
		logarithm_table[570] = 12'b000011_001010;
		logarithm_table[571] = 12'b000011_001010;
		logarithm_table[572] = 12'b000011_001010;
		logarithm_table[573] = 12'b000011_001010;
		logarithm_table[574] = 12'b000011_001011;
		logarithm_table[575] = 12'b000011_001011;
		logarithm_table[576] = 12'b000011_001011;
		logarithm_table[577] = 12'b000011_001011;
		logarithm_table[578] = 12'b000011_001011;
		logarithm_table[579] = 12'b000011_001011;
		logarithm_table[580] = 12'b000011_001100;
		logarithm_table[581] = 12'b000011_001100;
		logarithm_table[582] = 12'b000011_001100;
		logarithm_table[583] = 12'b000011_001100;
		logarithm_table[584] = 12'b000011_001100;
		logarithm_table[585] = 12'b000011_001100;
		logarithm_table[586] = 12'b000011_001100;
		logarithm_table[587] = 12'b000011_001101;
		logarithm_table[588] = 12'b000011_001101;
		logarithm_table[589] = 12'b000011_001101;
		logarithm_table[590] = 12'b000011_001101;
		logarithm_table[591] = 12'b000011_001101;
		logarithm_table[592] = 12'b000011_001101;
		logarithm_table[593] = 12'b000011_001110;
		logarithm_table[594] = 12'b000011_001110;
		logarithm_table[595] = 12'b000011_001110;
		logarithm_table[596] = 12'b000011_001110;
		logarithm_table[597] = 12'b000011_001110;
		logarithm_table[598] = 12'b000011_001110;
		logarithm_table[599] = 12'b000011_001110;
		logarithm_table[600] = 12'b000011_001111;
		logarithm_table[601] = 12'b000011_001111;
		logarithm_table[602] = 12'b000011_001111;
		logarithm_table[603] = 12'b000011_001111;
		logarithm_table[604] = 12'b000011_001111;
		logarithm_table[605] = 12'b000011_001111;
		logarithm_table[606] = 12'b000011_010000;
		logarithm_table[607] = 12'b000011_010000;
		logarithm_table[608] = 12'b000011_010000;
		logarithm_table[609] = 12'b000011_010000;
		logarithm_table[610] = 12'b000011_010000;
		logarithm_table[611] = 12'b000011_010000;
		logarithm_table[612] = 12'b000011_010000;
		logarithm_table[613] = 12'b000011_010001;
		logarithm_table[614] = 12'b000011_010001;
		logarithm_table[615] = 12'b000011_010001;
		logarithm_table[616] = 12'b000011_010001;
		logarithm_table[617] = 12'b000011_010001;
		logarithm_table[618] = 12'b000011_010001;
		logarithm_table[619] = 12'b000011_010010;
		logarithm_table[620] = 12'b000011_010010;
		logarithm_table[621] = 12'b000011_010010;
		logarithm_table[622] = 12'b000011_010010;
		logarithm_table[623] = 12'b000011_010010;
		logarithm_table[624] = 12'b000011_010010;
		logarithm_table[625] = 12'b000011_010010;
		logarithm_table[626] = 12'b000011_010011;
		logarithm_table[627] = 12'b000011_010011;
		logarithm_table[628] = 12'b000011_010011;
		logarithm_table[629] = 12'b000011_010011;
		logarithm_table[630] = 12'b000011_010011;
		logarithm_table[631] = 12'b000011_010011;
		logarithm_table[632] = 12'b000011_010011;
		logarithm_table[633] = 12'b000011_010100;
		logarithm_table[634] = 12'b000011_010100;
		logarithm_table[635] = 12'b000011_010100;
		logarithm_table[636] = 12'b000011_010100;
		logarithm_table[637] = 12'b000011_010100;
		logarithm_table[638] = 12'b000011_010100;
		logarithm_table[639] = 12'b000011_010100;
		logarithm_table[640] = 12'b000011_010101;
		logarithm_table[641] = 12'b000011_010101;
		logarithm_table[642] = 12'b000011_010101;
		logarithm_table[643] = 12'b000011_010101;
		logarithm_table[644] = 12'b000011_010101;
		logarithm_table[645] = 12'b000011_010101;
		logarithm_table[646] = 12'b000011_010101;
		logarithm_table[647] = 12'b000011_010110;
		logarithm_table[648] = 12'b000011_010110;
		logarithm_table[649] = 12'b000011_010110;
		logarithm_table[650] = 12'b000011_010110;
		logarithm_table[651] = 12'b000011_010110;
		logarithm_table[652] = 12'b000011_010110;
		logarithm_table[653] = 12'b000011_010110;
		logarithm_table[654] = 12'b000011_010111;
		logarithm_table[655] = 12'b000011_010111;
		logarithm_table[656] = 12'b000011_010111;
		logarithm_table[657] = 12'b000011_010111;
		logarithm_table[658] = 12'b000011_010111;
		logarithm_table[659] = 12'b000011_010111;
		logarithm_table[660] = 12'b000011_010111;
		logarithm_table[661] = 12'b000011_011000;
		logarithm_table[662] = 12'b000011_011000;
		logarithm_table[663] = 12'b000011_011000;
		logarithm_table[664] = 12'b000011_011000;
		logarithm_table[665] = 12'b000011_011000;
		logarithm_table[666] = 12'b000011_011000;
		logarithm_table[667] = 12'b000011_011000;
		logarithm_table[668] = 12'b000011_011001;
		logarithm_table[669] = 12'b000011_011001;
		logarithm_table[670] = 12'b000011_011001;
		logarithm_table[671] = 12'b000011_011001;
		logarithm_table[672] = 12'b000011_011001;
		logarithm_table[673] = 12'b000011_011001;
		logarithm_table[674] = 12'b000011_011001;
		logarithm_table[675] = 12'b000011_011010;
		logarithm_table[676] = 12'b000011_011010;
		logarithm_table[677] = 12'b000011_011010;
		logarithm_table[678] = 12'b000011_011010;
		logarithm_table[679] = 12'b000011_011010;
		logarithm_table[680] = 12'b000011_011010;
		logarithm_table[681] = 12'b000011_011010;
		logarithm_table[682] = 12'b000011_011010;
		logarithm_table[683] = 12'b000011_011011;
		logarithm_table[684] = 12'b000011_011011;
		logarithm_table[685] = 12'b000011_011011;
		logarithm_table[686] = 12'b000011_011011;
		logarithm_table[687] = 12'b000011_011011;
		logarithm_table[688] = 12'b000011_011011;
		logarithm_table[689] = 12'b000011_011011;
		logarithm_table[690] = 12'b000011_011100;
		logarithm_table[691] = 12'b000011_011100;
		logarithm_table[692] = 12'b000011_011100;
		logarithm_table[693] = 12'b000011_011100;
		logarithm_table[694] = 12'b000011_011100;
		logarithm_table[695] = 12'b000011_011100;
		logarithm_table[696] = 12'b000011_011100;
		logarithm_table[697] = 12'b000011_011100;
		logarithm_table[698] = 12'b000011_011101;
		logarithm_table[699] = 12'b000011_011101;
		logarithm_table[700] = 12'b000011_011101;
		logarithm_table[701] = 12'b000011_011101;
		logarithm_table[702] = 12'b000011_011101;
		logarithm_table[703] = 12'b000011_011101;
		logarithm_table[704] = 12'b000011_011101;
		logarithm_table[705] = 12'b000011_011110;
		logarithm_table[706] = 12'b000011_011110;
		logarithm_table[707] = 12'b000011_011110;
		logarithm_table[708] = 12'b000011_011110;
		logarithm_table[709] = 12'b000011_011110;
		logarithm_table[710] = 12'b000011_011110;
		logarithm_table[711] = 12'b000011_011110;
		logarithm_table[712] = 12'b000011_011110;
		logarithm_table[713] = 12'b000011_011111;
		logarithm_table[714] = 12'b000011_011111;
		logarithm_table[715] = 12'b000011_011111;
		logarithm_table[716] = 12'b000011_011111;
		logarithm_table[717] = 12'b000011_011111;
		logarithm_table[718] = 12'b000011_011111;
		logarithm_table[719] = 12'b000011_011111;
		logarithm_table[720] = 12'b000011_011111;
		logarithm_table[721] = 12'b000011_100000;
		logarithm_table[722] = 12'b000011_100000;
		logarithm_table[723] = 12'b000011_100000;
		logarithm_table[724] = 12'b000011_100000;
		logarithm_table[725] = 12'b000011_100000;
		logarithm_table[726] = 12'b000011_100000;
		logarithm_table[727] = 12'b000011_100000;
		logarithm_table[728] = 12'b000011_100000;
		logarithm_table[729] = 12'b000011_100001;
		logarithm_table[730] = 12'b000011_100001;
		logarithm_table[731] = 12'b000011_100001;
		logarithm_table[732] = 12'b000011_100001;
		logarithm_table[733] = 12'b000011_100001;
		logarithm_table[734] = 12'b000011_100001;
		logarithm_table[735] = 12'b000011_100001;
		logarithm_table[736] = 12'b000011_100010;
		logarithm_table[737] = 12'b000011_100010;
		logarithm_table[738] = 12'b000011_100010;
		logarithm_table[739] = 12'b000011_100010;
		logarithm_table[740] = 12'b000011_100010;
		logarithm_table[741] = 12'b000011_100010;
		logarithm_table[742] = 12'b000011_100010;
		logarithm_table[743] = 12'b000011_100010;
		logarithm_table[744] = 12'b000011_100011;
		logarithm_table[745] = 12'b000011_100011;
		logarithm_table[746] = 12'b000011_100011;
		logarithm_table[747] = 12'b000011_100011;
		logarithm_table[748] = 12'b000011_100011;
		logarithm_table[749] = 12'b000011_100011;
		logarithm_table[750] = 12'b000011_100011;
		logarithm_table[751] = 12'b000011_100011;
		logarithm_table[752] = 12'b000011_100011;
		logarithm_table[753] = 12'b000011_100100;
		logarithm_table[754] = 12'b000011_100100;
		logarithm_table[755] = 12'b000011_100100;
		logarithm_table[756] = 12'b000011_100100;
		logarithm_table[757] = 12'b000011_100100;
		logarithm_table[758] = 12'b000011_100100;
		logarithm_table[759] = 12'b000011_100100;
		logarithm_table[760] = 12'b000011_100100;
		logarithm_table[761] = 12'b000011_100101;
		logarithm_table[762] = 12'b000011_100101;
		logarithm_table[763] = 12'b000011_100101;
		logarithm_table[764] = 12'b000011_100101;
		logarithm_table[765] = 12'b000011_100101;
		logarithm_table[766] = 12'b000011_100101;
		logarithm_table[767] = 12'b000011_100101;
		logarithm_table[768] = 12'b000011_100101;
		logarithm_table[769] = 12'b000011_100110;
		logarithm_table[770] = 12'b000011_100110;
		logarithm_table[771] = 12'b000011_100110;
		logarithm_table[772] = 12'b000011_100110;
		logarithm_table[773] = 12'b000011_100110;
		logarithm_table[774] = 12'b000011_100110;
		logarithm_table[775] = 12'b000011_100110;
		logarithm_table[776] = 12'b000011_100110;
		logarithm_table[777] = 12'b000011_100111;
		logarithm_table[778] = 12'b000011_100111;
		logarithm_table[779] = 12'b000011_100111;
		logarithm_table[780] = 12'b000011_100111;
		logarithm_table[781] = 12'b000011_100111;
		logarithm_table[782] = 12'b000011_100111;
		logarithm_table[783] = 12'b000011_100111;
		logarithm_table[784] = 12'b000011_100111;
		logarithm_table[785] = 12'b000011_100111;
		logarithm_table[786] = 12'b000011_101000;
		logarithm_table[787] = 12'b000011_101000;
		logarithm_table[788] = 12'b000011_101000;
		logarithm_table[789] = 12'b000011_101000;
		logarithm_table[790] = 12'b000011_101000;
		logarithm_table[791] = 12'b000011_101000;
		logarithm_table[792] = 12'b000011_101000;
		logarithm_table[793] = 12'b000011_101000;
		logarithm_table[794] = 12'b000011_101001;
		logarithm_table[795] = 12'b000011_101001;
		logarithm_table[796] = 12'b000011_101001;
		logarithm_table[797] = 12'b000011_101001;
		logarithm_table[798] = 12'b000011_101001;
		logarithm_table[799] = 12'b000011_101001;
		logarithm_table[800] = 12'b000011_101001;
		logarithm_table[801] = 12'b000011_101001;
		logarithm_table[802] = 12'b000011_101001;
		logarithm_table[803] = 12'b000011_101010;
		logarithm_table[804] = 12'b000011_101010;
		logarithm_table[805] = 12'b000011_101010;
		logarithm_table[806] = 12'b000011_101010;
		logarithm_table[807] = 12'b000011_101010;
		logarithm_table[808] = 12'b000011_101010;
		logarithm_table[809] = 12'b000011_101010;
		logarithm_table[810] = 12'b000011_101010;
		logarithm_table[811] = 12'b000011_101010;
		logarithm_table[812] = 12'b000011_101011;
		logarithm_table[813] = 12'b000011_101011;
		logarithm_table[814] = 12'b000011_101011;
		logarithm_table[815] = 12'b000011_101011;
		logarithm_table[816] = 12'b000011_101011;
		logarithm_table[817] = 12'b000011_101011;
		logarithm_table[818] = 12'b000011_101011;
		logarithm_table[819] = 12'b000011_101011;
		logarithm_table[820] = 12'b000011_101011;
		logarithm_table[821] = 12'b000011_101100;
		logarithm_table[822] = 12'b000011_101100;
		logarithm_table[823] = 12'b000011_101100;
		logarithm_table[824] = 12'b000011_101100;
		logarithm_table[825] = 12'b000011_101100;
		logarithm_table[826] = 12'b000011_101100;
		logarithm_table[827] = 12'b000011_101100;
		logarithm_table[828] = 12'b000011_101100;
		logarithm_table[829] = 12'b000011_101100;
		logarithm_table[830] = 12'b000011_101101;
		logarithm_table[831] = 12'b000011_101101;
		logarithm_table[832] = 12'b000011_101101;
		logarithm_table[833] = 12'b000011_101101;
		logarithm_table[834] = 12'b000011_101101;
		logarithm_table[835] = 12'b000011_101101;
		logarithm_table[836] = 12'b000011_101101;
		logarithm_table[837] = 12'b000011_101101;
		logarithm_table[838] = 12'b000011_101101;
		logarithm_table[839] = 12'b000011_101110;
		logarithm_table[840] = 12'b000011_101110;
		logarithm_table[841] = 12'b000011_101110;
		logarithm_table[842] = 12'b000011_101110;
		logarithm_table[843] = 12'b000011_101110;
		logarithm_table[844] = 12'b000011_101110;
		logarithm_table[845] = 12'b000011_101110;
		logarithm_table[846] = 12'b000011_101110;
		logarithm_table[847] = 12'b000011_101110;
		logarithm_table[848] = 12'b000011_101111;
		logarithm_table[849] = 12'b000011_101111;
		logarithm_table[850] = 12'b000011_101111;
		logarithm_table[851] = 12'b000011_101111;
		logarithm_table[852] = 12'b000011_101111;
		logarithm_table[853] = 12'b000011_101111;
		logarithm_table[854] = 12'b000011_101111;
		logarithm_table[855] = 12'b000011_101111;
		logarithm_table[856] = 12'b000011_101111;
		logarithm_table[857] = 12'b000011_110000;
		logarithm_table[858] = 12'b000011_110000;
		logarithm_table[859] = 12'b000011_110000;
		logarithm_table[860] = 12'b000011_110000;
		logarithm_table[861] = 12'b000011_110000;
		logarithm_table[862] = 12'b000011_110000;
		logarithm_table[863] = 12'b000011_110000;
		logarithm_table[864] = 12'b000011_110000;
		logarithm_table[865] = 12'b000011_110000;
		logarithm_table[866] = 12'b000011_110001;
		logarithm_table[867] = 12'b000011_110001;
		logarithm_table[868] = 12'b000011_110001;
		logarithm_table[869] = 12'b000011_110001;
		logarithm_table[870] = 12'b000011_110001;
		logarithm_table[871] = 12'b000011_110001;
		logarithm_table[872] = 12'b000011_110001;
		logarithm_table[873] = 12'b000011_110001;
		logarithm_table[874] = 12'b000011_110001;
		logarithm_table[875] = 12'b000011_110001;
		logarithm_table[876] = 12'b000011_110010;
		logarithm_table[877] = 12'b000011_110010;
		logarithm_table[878] = 12'b000011_110010;
		logarithm_table[879] = 12'b000011_110010;
		logarithm_table[880] = 12'b000011_110010;
		logarithm_table[881] = 12'b000011_110010;
		logarithm_table[882] = 12'b000011_110010;
		logarithm_table[883] = 12'b000011_110010;
		logarithm_table[884] = 12'b000011_110010;
		logarithm_table[885] = 12'b000011_110011;
		logarithm_table[886] = 12'b000011_110011;
		logarithm_table[887] = 12'b000011_110011;
		logarithm_table[888] = 12'b000011_110011;
		logarithm_table[889] = 12'b000011_110011;
		logarithm_table[890] = 12'b000011_110011;
		logarithm_table[891] = 12'b000011_110011;
		logarithm_table[892] = 12'b000011_110011;
		logarithm_table[893] = 12'b000011_110011;
		logarithm_table[894] = 12'b000011_110011;
		logarithm_table[895] = 12'b000011_110100;
		logarithm_table[896] = 12'b000011_110100;
		logarithm_table[897] = 12'b000011_110100;
		logarithm_table[898] = 12'b000011_110100;
		logarithm_table[899] = 12'b000011_110100;
		logarithm_table[900] = 12'b000011_110100;
		logarithm_table[901] = 12'b000011_110100;
		logarithm_table[902] = 12'b000011_110100;
		logarithm_table[903] = 12'b000011_110100;
		logarithm_table[904] = 12'b000011_110100;
		logarithm_table[905] = 12'b000011_110101;
		logarithm_table[906] = 12'b000011_110101;
		logarithm_table[907] = 12'b000011_110101;
		logarithm_table[908] = 12'b000011_110101;
		logarithm_table[909] = 12'b000011_110101;
		logarithm_table[910] = 12'b000011_110101;
		logarithm_table[911] = 12'b000011_110101;
		logarithm_table[912] = 12'b000011_110101;
		logarithm_table[913] = 12'b000011_110101;
		logarithm_table[914] = 12'b000011_110110;
		logarithm_table[915] = 12'b000011_110110;
		logarithm_table[916] = 12'b000011_110110;
		logarithm_table[917] = 12'b000011_110110;
		logarithm_table[918] = 12'b000011_110110;
		logarithm_table[919] = 12'b000011_110110;
		logarithm_table[920] = 12'b000011_110110;
		logarithm_table[921] = 12'b000011_110110;
		logarithm_table[922] = 12'b000011_110110;
		logarithm_table[923] = 12'b000011_110110;
		logarithm_table[924] = 12'b000011_110111;
		logarithm_table[925] = 12'b000011_110111;
		logarithm_table[926] = 12'b000011_110111;
		logarithm_table[927] = 12'b000011_110111;
		logarithm_table[928] = 12'b000011_110111;
		logarithm_table[929] = 12'b000011_110111;
		logarithm_table[930] = 12'b000011_110111;
		logarithm_table[931] = 12'b000011_110111;
		logarithm_table[932] = 12'b000011_110111;
		logarithm_table[933] = 12'b000011_110111;
		logarithm_table[934] = 12'b000011_111000;
		logarithm_table[935] = 12'b000011_111000;
		logarithm_table[936] = 12'b000011_111000;
		logarithm_table[937] = 12'b000011_111000;
		logarithm_table[938] = 12'b000011_111000;
		logarithm_table[939] = 12'b000011_111000;
		logarithm_table[940] = 12'b000011_111000;
		logarithm_table[941] = 12'b000011_111000;
		logarithm_table[942] = 12'b000011_111000;
		logarithm_table[943] = 12'b000011_111000;
		logarithm_table[944] = 12'b000011_111000;
		logarithm_table[945] = 12'b000011_111001;
		logarithm_table[946] = 12'b000011_111001;
		logarithm_table[947] = 12'b000011_111001;
		logarithm_table[948] = 12'b000011_111001;
		logarithm_table[949] = 12'b000011_111001;
		logarithm_table[950] = 12'b000011_111001;
		logarithm_table[951] = 12'b000011_111001;
		logarithm_table[952] = 12'b000011_111001;
		logarithm_table[953] = 12'b000011_111001;
		logarithm_table[954] = 12'b000011_111001;
		logarithm_table[955] = 12'b000011_111010;
		logarithm_table[956] = 12'b000011_111010;
		logarithm_table[957] = 12'b000011_111010;
		logarithm_table[958] = 12'b000011_111010;
		logarithm_table[959] = 12'b000011_111010;
		logarithm_table[960] = 12'b000011_111010;
		logarithm_table[961] = 12'b000011_111010;
		logarithm_table[962] = 12'b000011_111010;
		logarithm_table[963] = 12'b000011_111010;
		logarithm_table[964] = 12'b000011_111010;
		logarithm_table[965] = 12'b000011_111011;
		logarithm_table[966] = 12'b000011_111011;
		logarithm_table[967] = 12'b000011_111011;
		logarithm_table[968] = 12'b000011_111011;
		logarithm_table[969] = 12'b000011_111011;
		logarithm_table[970] = 12'b000011_111011;
		logarithm_table[971] = 12'b000011_111011;
		logarithm_table[972] = 12'b000011_111011;
		logarithm_table[973] = 12'b000011_111011;
		logarithm_table[974] = 12'b000011_111011;
		logarithm_table[975] = 12'b000011_111011;
		logarithm_table[976] = 12'b000011_111100;
		logarithm_table[977] = 12'b000011_111100;
		logarithm_table[978] = 12'b000011_111100;
		logarithm_table[979] = 12'b000011_111100;
		logarithm_table[980] = 12'b000011_111100;
		logarithm_table[981] = 12'b000011_111100;
		logarithm_table[982] = 12'b000011_111100;
		logarithm_table[983] = 12'b000011_111100;
		logarithm_table[984] = 12'b000011_111100;
		logarithm_table[985] = 12'b000011_111100;
		logarithm_table[986] = 12'b000011_111101;
		logarithm_table[987] = 12'b000011_111101;
		logarithm_table[988] = 12'b000011_111101;
		logarithm_table[989] = 12'b000011_111101;
		logarithm_table[990] = 12'b000011_111101;
		logarithm_table[991] = 12'b000011_111101;
		logarithm_table[992] = 12'b000011_111101;
		logarithm_table[993] = 12'b000011_111101;
		logarithm_table[994] = 12'b000011_111101;
		logarithm_table[995] = 12'b000011_111101;
		logarithm_table[996] = 12'b000011_111101;
		logarithm_table[997] = 12'b000011_111110;
		logarithm_table[998] = 12'b000011_111110;
		logarithm_table[999] = 12'b000011_111110;
		logarithm_table[1000] = 12'b000011_111110;
		logarithm_table[1001] = 12'b000011_111110;
		logarithm_table[1002] = 12'b000011_111110;
		logarithm_table[1003] = 12'b000011_111110;
		logarithm_table[1004] = 12'b000011_111110;
		logarithm_table[1005] = 12'b000011_111110;
		logarithm_table[1006] = 12'b000011_111110;
		logarithm_table[1007] = 12'b000011_111110;
		logarithm_table[1008] = 12'b000011_111111;
		logarithm_table[1009] = 12'b000011_111111;
		logarithm_table[1010] = 12'b000011_111111;
		logarithm_table[1011] = 12'b000011_111111;
		logarithm_table[1012] = 12'b000011_111111;
		logarithm_table[1013] = 12'b000011_111111;
		logarithm_table[1014] = 12'b000011_111111;
		logarithm_table[1015] = 12'b000011_111111;
		logarithm_table[1016] = 12'b000011_111111;
		logarithm_table[1017] = 12'b000011_111111;
		logarithm_table[1018] = 12'b000011_111111;
		logarithm_table[1019] = 12'b000100_000000;
		logarithm_table[1020] = 12'b000100_000000;
		logarithm_table[1021] = 12'b000100_000000;
		logarithm_table[1022] = 12'b000100_000000;
		logarithm_table[1023] = 12'b000100_000000;
		logarithm_table[1024] = 12'b000100_000000;
		logarithm_table[1025] = 12'b000100_000000;
		logarithm_table[1026] = 12'b000100_000000;
		logarithm_table[1027] = 12'b000100_000000;
		logarithm_table[1028] = 12'b000100_000000;
		logarithm_table[1029] = 12'b000100_000000;
		logarithm_table[1030] = 12'b000100_000001;
		logarithm_table[1031] = 12'b000100_000001;
		logarithm_table[1032] = 12'b000100_000001;
		logarithm_table[1033] = 12'b000100_000001;
		logarithm_table[1034] = 12'b000100_000001;
		logarithm_table[1035] = 12'b000100_000001;
		logarithm_table[1036] = 12'b000100_000001;
		logarithm_table[1037] = 12'b000100_000001;
		logarithm_table[1038] = 12'b000100_000001;
		logarithm_table[1039] = 12'b000100_000001;
		logarithm_table[1040] = 12'b000100_000001;
		logarithm_table[1041] = 12'b000100_000010;
		logarithm_table[1042] = 12'b000100_000010;
		logarithm_table[1043] = 12'b000100_000010;
		logarithm_table[1044] = 12'b000100_000010;
		logarithm_table[1045] = 12'b000100_000010;
		logarithm_table[1046] = 12'b000100_000010;
		logarithm_table[1047] = 12'b000100_000010;
		logarithm_table[1048] = 12'b000100_000010;
		logarithm_table[1049] = 12'b000100_000010;
		logarithm_table[1050] = 12'b000100_000010;
		logarithm_table[1051] = 12'b000100_000010;
		logarithm_table[1052] = 12'b000100_000010;
		logarithm_table[1053] = 12'b000100_000011;
		logarithm_table[1054] = 12'b000100_000011;
		logarithm_table[1055] = 12'b000100_000011;
		logarithm_table[1056] = 12'b000100_000011;
		logarithm_table[1057] = 12'b000100_000011;
		logarithm_table[1058] = 12'b000100_000011;
		logarithm_table[1059] = 12'b000100_000011;
		logarithm_table[1060] = 12'b000100_000011;
		logarithm_table[1061] = 12'b000100_000011;
		logarithm_table[1062] = 12'b000100_000011;
		logarithm_table[1063] = 12'b000100_000011;
		logarithm_table[1064] = 12'b000100_000100;
		logarithm_table[1065] = 12'b000100_000100;
		logarithm_table[1066] = 12'b000100_000100;
		logarithm_table[1067] = 12'b000100_000100;
		logarithm_table[1068] = 12'b000100_000100;
		logarithm_table[1069] = 12'b000100_000100;
		logarithm_table[1070] = 12'b000100_000100;
		logarithm_table[1071] = 12'b000100_000100;
		logarithm_table[1072] = 12'b000100_000100;
		logarithm_table[1073] = 12'b000100_000100;
		logarithm_table[1074] = 12'b000100_000100;
		logarithm_table[1075] = 12'b000100_000100;
		logarithm_table[1076] = 12'b000100_000101;
		logarithm_table[1077] = 12'b000100_000101;
		logarithm_table[1078] = 12'b000100_000101;
		logarithm_table[1079] = 12'b000100_000101;
		logarithm_table[1080] = 12'b000100_000101;
		logarithm_table[1081] = 12'b000100_000101;
		logarithm_table[1082] = 12'b000100_000101;
		logarithm_table[1083] = 12'b000100_000101;
		logarithm_table[1084] = 12'b000100_000101;
		logarithm_table[1085] = 12'b000100_000101;
		logarithm_table[1086] = 12'b000100_000101;
		logarithm_table[1087] = 12'b000100_000110;
		logarithm_table[1088] = 12'b000100_000110;
		logarithm_table[1089] = 12'b000100_000110;
		logarithm_table[1090] = 12'b000100_000110;
		logarithm_table[1091] = 12'b000100_000110;
		logarithm_table[1092] = 12'b000100_000110;
		logarithm_table[1093] = 12'b000100_000110;
		logarithm_table[1094] = 12'b000100_000110;
		logarithm_table[1095] = 12'b000100_000110;
		logarithm_table[1096] = 12'b000100_000110;
		logarithm_table[1097] = 12'b000100_000110;
		logarithm_table[1098] = 12'b000100_000110;
		logarithm_table[1099] = 12'b000100_000111;
		logarithm_table[1100] = 12'b000100_000111;
		logarithm_table[1101] = 12'b000100_000111;
		logarithm_table[1102] = 12'b000100_000111;
		logarithm_table[1103] = 12'b000100_000111;
		logarithm_table[1104] = 12'b000100_000111;
		logarithm_table[1105] = 12'b000100_000111;
		logarithm_table[1106] = 12'b000100_000111;
		logarithm_table[1107] = 12'b000100_000111;
		logarithm_table[1108] = 12'b000100_000111;
		logarithm_table[1109] = 12'b000100_000111;
		logarithm_table[1110] = 12'b000100_000111;
		logarithm_table[1111] = 12'b000100_001000;
		logarithm_table[1112] = 12'b000100_001000;
		logarithm_table[1113] = 12'b000100_001000;
		logarithm_table[1114] = 12'b000100_001000;
		logarithm_table[1115] = 12'b000100_001000;
		logarithm_table[1116] = 12'b000100_001000;
		logarithm_table[1117] = 12'b000100_001000;
		logarithm_table[1118] = 12'b000100_001000;
		logarithm_table[1119] = 12'b000100_001000;
		logarithm_table[1120] = 12'b000100_001000;
		logarithm_table[1121] = 12'b000100_001000;
		logarithm_table[1122] = 12'b000100_001000;
		logarithm_table[1123] = 12'b000100_001001;
		logarithm_table[1124] = 12'b000100_001001;
		logarithm_table[1125] = 12'b000100_001001;
		logarithm_table[1126] = 12'b000100_001001;
		logarithm_table[1127] = 12'b000100_001001;
		logarithm_table[1128] = 12'b000100_001001;
		logarithm_table[1129] = 12'b000100_001001;
		logarithm_table[1130] = 12'b000100_001001;
		logarithm_table[1131] = 12'b000100_001001;
		logarithm_table[1132] = 12'b000100_001001;
		logarithm_table[1133] = 12'b000100_001001;
		logarithm_table[1134] = 12'b000100_001001;
		logarithm_table[1135] = 12'b000100_001010;
		logarithm_table[1136] = 12'b000100_001010;
		logarithm_table[1137] = 12'b000100_001010;
		logarithm_table[1138] = 12'b000100_001010;
		logarithm_table[1139] = 12'b000100_001010;
		logarithm_table[1140] = 12'b000100_001010;
		logarithm_table[1141] = 12'b000100_001010;
		logarithm_table[1142] = 12'b000100_001010;
		logarithm_table[1143] = 12'b000100_001010;
		logarithm_table[1144] = 12'b000100_001010;
		logarithm_table[1145] = 12'b000100_001010;
		logarithm_table[1146] = 12'b000100_001010;
		logarithm_table[1147] = 12'b000100_001010;
		logarithm_table[1148] = 12'b000100_001011;
		logarithm_table[1149] = 12'b000100_001011;
		logarithm_table[1150] = 12'b000100_001011;
		logarithm_table[1151] = 12'b000100_001011;
		logarithm_table[1152] = 12'b000100_001011;
		logarithm_table[1153] = 12'b000100_001011;
		logarithm_table[1154] = 12'b000100_001011;
		logarithm_table[1155] = 12'b000100_001011;
		logarithm_table[1156] = 12'b000100_001011;
		logarithm_table[1157] = 12'b000100_001011;
		logarithm_table[1158] = 12'b000100_001011;
		logarithm_table[1159] = 12'b000100_001011;
		logarithm_table[1160] = 12'b000100_001100;
		logarithm_table[1161] = 12'b000100_001100;
		logarithm_table[1162] = 12'b000100_001100;
		logarithm_table[1163] = 12'b000100_001100;
		logarithm_table[1164] = 12'b000100_001100;
		logarithm_table[1165] = 12'b000100_001100;
		logarithm_table[1166] = 12'b000100_001100;
		logarithm_table[1167] = 12'b000100_001100;
		logarithm_table[1168] = 12'b000100_001100;
		logarithm_table[1169] = 12'b000100_001100;
		logarithm_table[1170] = 12'b000100_001100;
		logarithm_table[1171] = 12'b000100_001100;
		logarithm_table[1172] = 12'b000100_001100;
		logarithm_table[1173] = 12'b000100_001101;
		logarithm_table[1174] = 12'b000100_001101;
		logarithm_table[1175] = 12'b000100_001101;
		logarithm_table[1176] = 12'b000100_001101;
		logarithm_table[1177] = 12'b000100_001101;
		logarithm_table[1178] = 12'b000100_001101;
		logarithm_table[1179] = 12'b000100_001101;
		logarithm_table[1180] = 12'b000100_001101;
		logarithm_table[1181] = 12'b000100_001101;
		logarithm_table[1182] = 12'b000100_001101;
		logarithm_table[1183] = 12'b000100_001101;
		logarithm_table[1184] = 12'b000100_001101;
		logarithm_table[1185] = 12'b000100_001101;
		logarithm_table[1186] = 12'b000100_001110;
		logarithm_table[1187] = 12'b000100_001110;
		logarithm_table[1188] = 12'b000100_001110;
		logarithm_table[1189] = 12'b000100_001110;
		logarithm_table[1190] = 12'b000100_001110;
		logarithm_table[1191] = 12'b000100_001110;
		logarithm_table[1192] = 12'b000100_001110;
		logarithm_table[1193] = 12'b000100_001110;
		logarithm_table[1194] = 12'b000100_001110;
		logarithm_table[1195] = 12'b000100_001110;
		logarithm_table[1196] = 12'b000100_001110;
		logarithm_table[1197] = 12'b000100_001110;
		logarithm_table[1198] = 12'b000100_001110;
		logarithm_table[1199] = 12'b000100_001111;
		logarithm_table[1200] = 12'b000100_001111;
		logarithm_table[1201] = 12'b000100_001111;
		logarithm_table[1202] = 12'b000100_001111;
		logarithm_table[1203] = 12'b000100_001111;
		logarithm_table[1204] = 12'b000100_001111;
		logarithm_table[1205] = 12'b000100_001111;
		logarithm_table[1206] = 12'b000100_001111;
		logarithm_table[1207] = 12'b000100_001111;
		logarithm_table[1208] = 12'b000100_001111;
		logarithm_table[1209] = 12'b000100_001111;
		logarithm_table[1210] = 12'b000100_001111;
		logarithm_table[1211] = 12'b000100_001111;
		logarithm_table[1212] = 12'b000100_010000;
		logarithm_table[1213] = 12'b000100_010000;
		logarithm_table[1214] = 12'b000100_010000;
		logarithm_table[1215] = 12'b000100_010000;
		logarithm_table[1216] = 12'b000100_010000;
		logarithm_table[1217] = 12'b000100_010000;
		logarithm_table[1218] = 12'b000100_010000;
		logarithm_table[1219] = 12'b000100_010000;
		logarithm_table[1220] = 12'b000100_010000;
		logarithm_table[1221] = 12'b000100_010000;
		logarithm_table[1222] = 12'b000100_010000;
		logarithm_table[1223] = 12'b000100_010000;
		logarithm_table[1224] = 12'b000100_010000;
		logarithm_table[1225] = 12'b000100_010001;
		logarithm_table[1226] = 12'b000100_010001;
		logarithm_table[1227] = 12'b000100_010001;
		logarithm_table[1228] = 12'b000100_010001;
		logarithm_table[1229] = 12'b000100_010001;
		logarithm_table[1230] = 12'b000100_010001;
		logarithm_table[1231] = 12'b000100_010001;
		logarithm_table[1232] = 12'b000100_010001;
		logarithm_table[1233] = 12'b000100_010001;
		logarithm_table[1234] = 12'b000100_010001;
		logarithm_table[1235] = 12'b000100_010001;
		logarithm_table[1236] = 12'b000100_010001;
		logarithm_table[1237] = 12'b000100_010001;
		logarithm_table[1238] = 12'b000100_010010;
		logarithm_table[1239] = 12'b000100_010010;
		logarithm_table[1240] = 12'b000100_010010;
		logarithm_table[1241] = 12'b000100_010010;
		logarithm_table[1242] = 12'b000100_010010;
		logarithm_table[1243] = 12'b000100_010010;
		logarithm_table[1244] = 12'b000100_010010;
		logarithm_table[1245] = 12'b000100_010010;
		logarithm_table[1246] = 12'b000100_010010;
		logarithm_table[1247] = 12'b000100_010010;
		logarithm_table[1248] = 12'b000100_010010;
		logarithm_table[1249] = 12'b000100_010010;
		logarithm_table[1250] = 12'b000100_010010;
		logarithm_table[1251] = 12'b000100_010010;
		logarithm_table[1252] = 12'b000100_010011;
		logarithm_table[1253] = 12'b000100_010011;
		logarithm_table[1254] = 12'b000100_010011;
		logarithm_table[1255] = 12'b000100_010011;
		logarithm_table[1256] = 12'b000100_010011;
		logarithm_table[1257] = 12'b000100_010011;
		logarithm_table[1258] = 12'b000100_010011;
		logarithm_table[1259] = 12'b000100_010011;
		logarithm_table[1260] = 12'b000100_010011;
		logarithm_table[1261] = 12'b000100_010011;
		logarithm_table[1262] = 12'b000100_010011;
		logarithm_table[1263] = 12'b000100_010011;
		logarithm_table[1264] = 12'b000100_010011;
		logarithm_table[1265] = 12'b000100_010100;
		logarithm_table[1266] = 12'b000100_010100;
		logarithm_table[1267] = 12'b000100_010100;
		logarithm_table[1268] = 12'b000100_010100;
		logarithm_table[1269] = 12'b000100_010100;
		logarithm_table[1270] = 12'b000100_010100;
		logarithm_table[1271] = 12'b000100_010100;
		logarithm_table[1272] = 12'b000100_010100;
		logarithm_table[1273] = 12'b000100_010100;
		logarithm_table[1274] = 12'b000100_010100;
		logarithm_table[1275] = 12'b000100_010100;
		logarithm_table[1276] = 12'b000100_010100;
		logarithm_table[1277] = 12'b000100_010100;
		logarithm_table[1278] = 12'b000100_010100;
		logarithm_table[1279] = 12'b000100_010101;
		logarithm_table[1280] = 12'b000100_010101;
		logarithm_table[1281] = 12'b000100_010101;
		logarithm_table[1282] = 12'b000100_010101;
		logarithm_table[1283] = 12'b000100_010101;
		logarithm_table[1284] = 12'b000100_010101;
		logarithm_table[1285] = 12'b000100_010101;
		logarithm_table[1286] = 12'b000100_010101;
		logarithm_table[1287] = 12'b000100_010101;
		logarithm_table[1288] = 12'b000100_010101;
		logarithm_table[1289] = 12'b000100_010101;
		logarithm_table[1290] = 12'b000100_010101;
		logarithm_table[1291] = 12'b000100_010101;
		logarithm_table[1292] = 12'b000100_010101;
		logarithm_table[1293] = 12'b000100_010110;
		logarithm_table[1294] = 12'b000100_010110;
		logarithm_table[1295] = 12'b000100_010110;
		logarithm_table[1296] = 12'b000100_010110;
		logarithm_table[1297] = 12'b000100_010110;
		logarithm_table[1298] = 12'b000100_010110;
		logarithm_table[1299] = 12'b000100_010110;
		logarithm_table[1300] = 12'b000100_010110;
		logarithm_table[1301] = 12'b000100_010110;
		logarithm_table[1302] = 12'b000100_010110;
		logarithm_table[1303] = 12'b000100_010110;
		logarithm_table[1304] = 12'b000100_010110;
		logarithm_table[1305] = 12'b000100_010110;
		logarithm_table[1306] = 12'b000100_010110;
		logarithm_table[1307] = 12'b000100_010111;
		logarithm_table[1308] = 12'b000100_010111;
		logarithm_table[1309] = 12'b000100_010111;
		logarithm_table[1310] = 12'b000100_010111;
		logarithm_table[1311] = 12'b000100_010111;
		logarithm_table[1312] = 12'b000100_010111;
		logarithm_table[1313] = 12'b000100_010111;
		logarithm_table[1314] = 12'b000100_010111;
		logarithm_table[1315] = 12'b000100_010111;
		logarithm_table[1316] = 12'b000100_010111;
		logarithm_table[1317] = 12'b000100_010111;
		logarithm_table[1318] = 12'b000100_010111;
		logarithm_table[1319] = 12'b000100_010111;
		logarithm_table[1320] = 12'b000100_010111;
		logarithm_table[1321] = 12'b000100_011000;
		logarithm_table[1322] = 12'b000100_011000;
		logarithm_table[1323] = 12'b000100_011000;
		logarithm_table[1324] = 12'b000100_011000;
		logarithm_table[1325] = 12'b000100_011000;
		logarithm_table[1326] = 12'b000100_011000;
		logarithm_table[1327] = 12'b000100_011000;
		logarithm_table[1328] = 12'b000100_011000;
		logarithm_table[1329] = 12'b000100_011000;
		logarithm_table[1330] = 12'b000100_011000;
		logarithm_table[1331] = 12'b000100_011000;
		logarithm_table[1332] = 12'b000100_011000;
		logarithm_table[1333] = 12'b000100_011000;
		logarithm_table[1334] = 12'b000100_011000;
		logarithm_table[1335] = 12'b000100_011000;
		logarithm_table[1336] = 12'b000100_011001;
		logarithm_table[1337] = 12'b000100_011001;
		logarithm_table[1338] = 12'b000100_011001;
		logarithm_table[1339] = 12'b000100_011001;
		logarithm_table[1340] = 12'b000100_011001;
		logarithm_table[1341] = 12'b000100_011001;
		logarithm_table[1342] = 12'b000100_011001;
		logarithm_table[1343] = 12'b000100_011001;
		logarithm_table[1344] = 12'b000100_011001;
		logarithm_table[1345] = 12'b000100_011001;
		logarithm_table[1346] = 12'b000100_011001;
		logarithm_table[1347] = 12'b000100_011001;
		logarithm_table[1348] = 12'b000100_011001;
		logarithm_table[1349] = 12'b000100_011001;
		logarithm_table[1350] = 12'b000100_011010;
		logarithm_table[1351] = 12'b000100_011010;
		logarithm_table[1352] = 12'b000100_011010;
		logarithm_table[1353] = 12'b000100_011010;
		logarithm_table[1354] = 12'b000100_011010;
		logarithm_table[1355] = 12'b000100_011010;
		logarithm_table[1356] = 12'b000100_011010;
		logarithm_table[1357] = 12'b000100_011010;
		logarithm_table[1358] = 12'b000100_011010;
		logarithm_table[1359] = 12'b000100_011010;
		logarithm_table[1360] = 12'b000100_011010;
		logarithm_table[1361] = 12'b000100_011010;
		logarithm_table[1362] = 12'b000100_011010;
		logarithm_table[1363] = 12'b000100_011010;
		logarithm_table[1364] = 12'b000100_011010;
		logarithm_table[1365] = 12'b000100_011011;
		logarithm_table[1366] = 12'b000100_011011;
		logarithm_table[1367] = 12'b000100_011011;
		logarithm_table[1368] = 12'b000100_011011;
		logarithm_table[1369] = 12'b000100_011011;
		logarithm_table[1370] = 12'b000100_011011;
		logarithm_table[1371] = 12'b000100_011011;
		logarithm_table[1372] = 12'b000100_011011;
		logarithm_table[1373] = 12'b000100_011011;
		logarithm_table[1374] = 12'b000100_011011;
		logarithm_table[1375] = 12'b000100_011011;
		logarithm_table[1376] = 12'b000100_011011;
		logarithm_table[1377] = 12'b000100_011011;
		logarithm_table[1378] = 12'b000100_011011;
		logarithm_table[1379] = 12'b000100_011011;
		logarithm_table[1380] = 12'b000100_011100;
		logarithm_table[1381] = 12'b000100_011100;
		logarithm_table[1382] = 12'b000100_011100;
		logarithm_table[1383] = 12'b000100_011100;
		logarithm_table[1384] = 12'b000100_011100;
		logarithm_table[1385] = 12'b000100_011100;
		logarithm_table[1386] = 12'b000100_011100;
		logarithm_table[1387] = 12'b000100_011100;
		logarithm_table[1388] = 12'b000100_011100;
		logarithm_table[1389] = 12'b000100_011100;
		logarithm_table[1390] = 12'b000100_011100;
		logarithm_table[1391] = 12'b000100_011100;
		logarithm_table[1392] = 12'b000100_011100;
		logarithm_table[1393] = 12'b000100_011100;
		logarithm_table[1394] = 12'b000100_011100;
		logarithm_table[1395] = 12'b000100_011101;
		logarithm_table[1396] = 12'b000100_011101;
		logarithm_table[1397] = 12'b000100_011101;
		logarithm_table[1398] = 12'b000100_011101;
		logarithm_table[1399] = 12'b000100_011101;
		logarithm_table[1400] = 12'b000100_011101;
		logarithm_table[1401] = 12'b000100_011101;
		logarithm_table[1402] = 12'b000100_011101;
		logarithm_table[1403] = 12'b000100_011101;
		logarithm_table[1404] = 12'b000100_011101;
		logarithm_table[1405] = 12'b000100_011101;
		logarithm_table[1406] = 12'b000100_011101;
		logarithm_table[1407] = 12'b000100_011101;
		logarithm_table[1408] = 12'b000100_011101;
		logarithm_table[1409] = 12'b000100_011101;
		logarithm_table[1410] = 12'b000100_011110;
		logarithm_table[1411] = 12'b000100_011110;
		logarithm_table[1412] = 12'b000100_011110;
		logarithm_table[1413] = 12'b000100_011110;
		logarithm_table[1414] = 12'b000100_011110;
		logarithm_table[1415] = 12'b000100_011110;
		logarithm_table[1416] = 12'b000100_011110;
		logarithm_table[1417] = 12'b000100_011110;
		logarithm_table[1418] = 12'b000100_011110;
		logarithm_table[1419] = 12'b000100_011110;
		logarithm_table[1420] = 12'b000100_011110;
		logarithm_table[1421] = 12'b000100_011110;
		logarithm_table[1422] = 12'b000100_011110;
		logarithm_table[1423] = 12'b000100_011110;
		logarithm_table[1424] = 12'b000100_011110;
		logarithm_table[1425] = 12'b000100_011111;
		logarithm_table[1426] = 12'b000100_011111;
		logarithm_table[1427] = 12'b000100_011111;
		logarithm_table[1428] = 12'b000100_011111;
		logarithm_table[1429] = 12'b000100_011111;
		logarithm_table[1430] = 12'b000100_011111;
		logarithm_table[1431] = 12'b000100_011111;
		logarithm_table[1432] = 12'b000100_011111;
		logarithm_table[1433] = 12'b000100_011111;
		logarithm_table[1434] = 12'b000100_011111;
		logarithm_table[1435] = 12'b000100_011111;
		logarithm_table[1436] = 12'b000100_011111;
		logarithm_table[1437] = 12'b000100_011111;
		logarithm_table[1438] = 12'b000100_011111;
		logarithm_table[1439] = 12'b000100_011111;
		logarithm_table[1440] = 12'b000100_011111;
		logarithm_table[1441] = 12'b000100_100000;
		logarithm_table[1442] = 12'b000100_100000;
		logarithm_table[1443] = 12'b000100_100000;
		logarithm_table[1444] = 12'b000100_100000;
		logarithm_table[1445] = 12'b000100_100000;
		logarithm_table[1446] = 12'b000100_100000;
		logarithm_table[1447] = 12'b000100_100000;
		logarithm_table[1448] = 12'b000100_100000;
		logarithm_table[1449] = 12'b000100_100000;
		logarithm_table[1450] = 12'b000100_100000;
		logarithm_table[1451] = 12'b000100_100000;
		logarithm_table[1452] = 12'b000100_100000;
		logarithm_table[1453] = 12'b000100_100000;
		logarithm_table[1454] = 12'b000100_100000;
		logarithm_table[1455] = 12'b000100_100000;
		logarithm_table[1456] = 12'b000100_100000;
		logarithm_table[1457] = 12'b000100_100001;
		logarithm_table[1458] = 12'b000100_100001;
		logarithm_table[1459] = 12'b000100_100001;
		logarithm_table[1460] = 12'b000100_100001;
		logarithm_table[1461] = 12'b000100_100001;
		logarithm_table[1462] = 12'b000100_100001;
		logarithm_table[1463] = 12'b000100_100001;
		logarithm_table[1464] = 12'b000100_100001;
		logarithm_table[1465] = 12'b000100_100001;
		logarithm_table[1466] = 12'b000100_100001;
		logarithm_table[1467] = 12'b000100_100001;
		logarithm_table[1468] = 12'b000100_100001;
		logarithm_table[1469] = 12'b000100_100001;
		logarithm_table[1470] = 12'b000100_100001;
		logarithm_table[1471] = 12'b000100_100001;
		logarithm_table[1472] = 12'b000100_100010;
		logarithm_table[1473] = 12'b000100_100010;
		logarithm_table[1474] = 12'b000100_100010;
		logarithm_table[1475] = 12'b000100_100010;
		logarithm_table[1476] = 12'b000100_100010;
		logarithm_table[1477] = 12'b000100_100010;
		logarithm_table[1478] = 12'b000100_100010;
		logarithm_table[1479] = 12'b000100_100010;
		logarithm_table[1480] = 12'b000100_100010;
		logarithm_table[1481] = 12'b000100_100010;
		logarithm_table[1482] = 12'b000100_100010;
		logarithm_table[1483] = 12'b000100_100010;
		logarithm_table[1484] = 12'b000100_100010;
		logarithm_table[1485] = 12'b000100_100010;
		logarithm_table[1486] = 12'b000100_100010;
		logarithm_table[1487] = 12'b000100_100010;
		logarithm_table[1488] = 12'b000100_100011;
		logarithm_table[1489] = 12'b000100_100011;
		logarithm_table[1490] = 12'b000100_100011;
		logarithm_table[1491] = 12'b000100_100011;
		logarithm_table[1492] = 12'b000100_100011;
		logarithm_table[1493] = 12'b000100_100011;
		logarithm_table[1494] = 12'b000100_100011;
		logarithm_table[1495] = 12'b000100_100011;
		logarithm_table[1496] = 12'b000100_100011;
		logarithm_table[1497] = 12'b000100_100011;
		logarithm_table[1498] = 12'b000100_100011;
		logarithm_table[1499] = 12'b000100_100011;
		logarithm_table[1500] = 12'b000100_100011;
		logarithm_table[1501] = 12'b000100_100011;
		logarithm_table[1502] = 12'b000100_100011;
		logarithm_table[1503] = 12'b000100_100011;
		logarithm_table[1504] = 12'b000100_100011;
		logarithm_table[1505] = 12'b000100_100100;
		logarithm_table[1506] = 12'b000100_100100;
		logarithm_table[1507] = 12'b000100_100100;
		logarithm_table[1508] = 12'b000100_100100;
		logarithm_table[1509] = 12'b000100_100100;
		logarithm_table[1510] = 12'b000100_100100;
		logarithm_table[1511] = 12'b000100_100100;
		logarithm_table[1512] = 12'b000100_100100;
		logarithm_table[1513] = 12'b000100_100100;
		logarithm_table[1514] = 12'b000100_100100;
		logarithm_table[1515] = 12'b000100_100100;
		logarithm_table[1516] = 12'b000100_100100;
		logarithm_table[1517] = 12'b000100_100100;
		logarithm_table[1518] = 12'b000100_100100;
		logarithm_table[1519] = 12'b000100_100100;
		logarithm_table[1520] = 12'b000100_100100;
		logarithm_table[1521] = 12'b000100_100101;
		logarithm_table[1522] = 12'b000100_100101;
		logarithm_table[1523] = 12'b000100_100101;
		logarithm_table[1524] = 12'b000100_100101;
		logarithm_table[1525] = 12'b000100_100101;
		logarithm_table[1526] = 12'b000100_100101;
		logarithm_table[1527] = 12'b000100_100101;
		logarithm_table[1528] = 12'b000100_100101;
		logarithm_table[1529] = 12'b000100_100101;
		logarithm_table[1530] = 12'b000100_100101;
		logarithm_table[1531] = 12'b000100_100101;
		logarithm_table[1532] = 12'b000100_100101;
		logarithm_table[1533] = 12'b000100_100101;
		logarithm_table[1534] = 12'b000100_100101;
		logarithm_table[1535] = 12'b000100_100101;
		logarithm_table[1536] = 12'b000100_100101;
		logarithm_table[1537] = 12'b000100_100101;
		logarithm_table[1538] = 12'b000100_100110;
		logarithm_table[1539] = 12'b000100_100110;
		logarithm_table[1540] = 12'b000100_100110;
		logarithm_table[1541] = 12'b000100_100110;
		logarithm_table[1542] = 12'b000100_100110;
		logarithm_table[1543] = 12'b000100_100110;
		logarithm_table[1544] = 12'b000100_100110;
		logarithm_table[1545] = 12'b000100_100110;
		logarithm_table[1546] = 12'b000100_100110;
		logarithm_table[1547] = 12'b000100_100110;
		logarithm_table[1548] = 12'b000100_100110;
		logarithm_table[1549] = 12'b000100_100110;
		logarithm_table[1550] = 12'b000100_100110;
		logarithm_table[1551] = 12'b000100_100110;
		logarithm_table[1552] = 12'b000100_100110;
		logarithm_table[1553] = 12'b000100_100110;
		logarithm_table[1554] = 12'b000100_100111;
		logarithm_table[1555] = 12'b000100_100111;
		logarithm_table[1556] = 12'b000100_100111;
		logarithm_table[1557] = 12'b000100_100111;
		logarithm_table[1558] = 12'b000100_100111;
		logarithm_table[1559] = 12'b000100_100111;
		logarithm_table[1560] = 12'b000100_100111;
		logarithm_table[1561] = 12'b000100_100111;
		logarithm_table[1562] = 12'b000100_100111;
		logarithm_table[1563] = 12'b000100_100111;
		logarithm_table[1564] = 12'b000100_100111;
		logarithm_table[1565] = 12'b000100_100111;
		logarithm_table[1566] = 12'b000100_100111;
		logarithm_table[1567] = 12'b000100_100111;
		logarithm_table[1568] = 12'b000100_100111;
		logarithm_table[1569] = 12'b000100_100111;
		logarithm_table[1570] = 12'b000100_100111;
		logarithm_table[1571] = 12'b000100_101000;
		logarithm_table[1572] = 12'b000100_101000;
		logarithm_table[1573] = 12'b000100_101000;
		logarithm_table[1574] = 12'b000100_101000;
		logarithm_table[1575] = 12'b000100_101000;
		logarithm_table[1576] = 12'b000100_101000;
		logarithm_table[1577] = 12'b000100_101000;
		logarithm_table[1578] = 12'b000100_101000;
		logarithm_table[1579] = 12'b000100_101000;
		logarithm_table[1580] = 12'b000100_101000;
		logarithm_table[1581] = 12'b000100_101000;
		logarithm_table[1582] = 12'b000100_101000;
		logarithm_table[1583] = 12'b000100_101000;
		logarithm_table[1584] = 12'b000100_101000;
		logarithm_table[1585] = 12'b000100_101000;
		logarithm_table[1586] = 12'b000100_101000;
		logarithm_table[1587] = 12'b000100_101000;
		logarithm_table[1588] = 12'b000100_101001;
		logarithm_table[1589] = 12'b000100_101001;
		logarithm_table[1590] = 12'b000100_101001;
		logarithm_table[1591] = 12'b000100_101001;
		logarithm_table[1592] = 12'b000100_101001;
		logarithm_table[1593] = 12'b000100_101001;
		logarithm_table[1594] = 12'b000100_101001;
		logarithm_table[1595] = 12'b000100_101001;
		logarithm_table[1596] = 12'b000100_101001;
		logarithm_table[1597] = 12'b000100_101001;
		logarithm_table[1598] = 12'b000100_101001;
		logarithm_table[1599] = 12'b000100_101001;
		logarithm_table[1600] = 12'b000100_101001;
		logarithm_table[1601] = 12'b000100_101001;
		logarithm_table[1602] = 12'b000100_101001;
		logarithm_table[1603] = 12'b000100_101001;
		logarithm_table[1604] = 12'b000100_101001;
		logarithm_table[1605] = 12'b000100_101001;
		logarithm_table[1606] = 12'b000100_101010;
		logarithm_table[1607] = 12'b000100_101010;
		logarithm_table[1608] = 12'b000100_101010;
		logarithm_table[1609] = 12'b000100_101010;
		logarithm_table[1610] = 12'b000100_101010;
		logarithm_table[1611] = 12'b000100_101010;
		logarithm_table[1612] = 12'b000100_101010;
		logarithm_table[1613] = 12'b000100_101010;
		logarithm_table[1614] = 12'b000100_101010;
		logarithm_table[1615] = 12'b000100_101010;
		logarithm_table[1616] = 12'b000100_101010;
		logarithm_table[1617] = 12'b000100_101010;
		logarithm_table[1618] = 12'b000100_101010;
		logarithm_table[1619] = 12'b000100_101010;
		logarithm_table[1620] = 12'b000100_101010;
		logarithm_table[1621] = 12'b000100_101010;
		logarithm_table[1622] = 12'b000100_101010;
		logarithm_table[1623] = 12'b000100_101011;
		logarithm_table[1624] = 12'b000100_101011;
		logarithm_table[1625] = 12'b000100_101011;
		logarithm_table[1626] = 12'b000100_101011;
		logarithm_table[1627] = 12'b000100_101011;
		logarithm_table[1628] = 12'b000100_101011;
		logarithm_table[1629] = 12'b000100_101011;
		logarithm_table[1630] = 12'b000100_101011;
		logarithm_table[1631] = 12'b000100_101011;
		logarithm_table[1632] = 12'b000100_101011;
		logarithm_table[1633] = 12'b000100_101011;
		logarithm_table[1634] = 12'b000100_101011;
		logarithm_table[1635] = 12'b000100_101011;
		logarithm_table[1636] = 12'b000100_101011;
		logarithm_table[1637] = 12'b000100_101011;
		logarithm_table[1638] = 12'b000100_101011;
		logarithm_table[1639] = 12'b000100_101011;
		logarithm_table[1640] = 12'b000100_101011;
		logarithm_table[1641] = 12'b000100_101100;
		logarithm_table[1642] = 12'b000100_101100;
		logarithm_table[1643] = 12'b000100_101100;
		logarithm_table[1644] = 12'b000100_101100;
		logarithm_table[1645] = 12'b000100_101100;
		logarithm_table[1646] = 12'b000100_101100;
		logarithm_table[1647] = 12'b000100_101100;
		logarithm_table[1648] = 12'b000100_101100;
		logarithm_table[1649] = 12'b000100_101100;
		logarithm_table[1650] = 12'b000100_101100;
		logarithm_table[1651] = 12'b000100_101100;
		logarithm_table[1652] = 12'b000100_101100;
		logarithm_table[1653] = 12'b000100_101100;
		logarithm_table[1654] = 12'b000100_101100;
		logarithm_table[1655] = 12'b000100_101100;
		logarithm_table[1656] = 12'b000100_101100;
		logarithm_table[1657] = 12'b000100_101100;
		logarithm_table[1658] = 12'b000100_101100;
		logarithm_table[1659] = 12'b000100_101101;
		logarithm_table[1660] = 12'b000100_101101;
		logarithm_table[1661] = 12'b000100_101101;
		logarithm_table[1662] = 12'b000100_101101;
		logarithm_table[1663] = 12'b000100_101101;
		logarithm_table[1664] = 12'b000100_101101;
		logarithm_table[1665] = 12'b000100_101101;
		logarithm_table[1666] = 12'b000100_101101;
		logarithm_table[1667] = 12'b000100_101101;
		logarithm_table[1668] = 12'b000100_101101;
		logarithm_table[1669] = 12'b000100_101101;
		logarithm_table[1670] = 12'b000100_101101;
		logarithm_table[1671] = 12'b000100_101101;
		logarithm_table[1672] = 12'b000100_101101;
		logarithm_table[1673] = 12'b000100_101101;
		logarithm_table[1674] = 12'b000100_101101;
		logarithm_table[1675] = 12'b000100_101101;
		logarithm_table[1676] = 12'b000100_101101;
		logarithm_table[1677] = 12'b000100_101110;
		logarithm_table[1678] = 12'b000100_101110;
		logarithm_table[1679] = 12'b000100_101110;
		logarithm_table[1680] = 12'b000100_101110;
		logarithm_table[1681] = 12'b000100_101110;
		logarithm_table[1682] = 12'b000100_101110;
		logarithm_table[1683] = 12'b000100_101110;
		logarithm_table[1684] = 12'b000100_101110;
		logarithm_table[1685] = 12'b000100_101110;
		logarithm_table[1686] = 12'b000100_101110;
		logarithm_table[1687] = 12'b000100_101110;
		logarithm_table[1688] = 12'b000100_101110;
		logarithm_table[1689] = 12'b000100_101110;
		logarithm_table[1690] = 12'b000100_101110;
		logarithm_table[1691] = 12'b000100_101110;
		logarithm_table[1692] = 12'b000100_101110;
		logarithm_table[1693] = 12'b000100_101110;
		logarithm_table[1694] = 12'b000100_101110;
		logarithm_table[1695] = 12'b000100_101111;
		logarithm_table[1696] = 12'b000100_101111;
		logarithm_table[1697] = 12'b000100_101111;
		logarithm_table[1698] = 12'b000100_101111;
		logarithm_table[1699] = 12'b000100_101111;
		logarithm_table[1700] = 12'b000100_101111;
		logarithm_table[1701] = 12'b000100_101111;
		logarithm_table[1702] = 12'b000100_101111;
		logarithm_table[1703] = 12'b000100_101111;
		logarithm_table[1704] = 12'b000100_101111;
		logarithm_table[1705] = 12'b000100_101111;
		logarithm_table[1706] = 12'b000100_101111;
		logarithm_table[1707] = 12'b000100_101111;
		logarithm_table[1708] = 12'b000100_101111;
		logarithm_table[1709] = 12'b000100_101111;
		logarithm_table[1710] = 12'b000100_101111;
		logarithm_table[1711] = 12'b000100_101111;
		logarithm_table[1712] = 12'b000100_101111;
		logarithm_table[1713] = 12'b000100_110000;
		logarithm_table[1714] = 12'b000100_110000;
		logarithm_table[1715] = 12'b000100_110000;
		logarithm_table[1716] = 12'b000100_110000;
		logarithm_table[1717] = 12'b000100_110000;
		logarithm_table[1718] = 12'b000100_110000;
		logarithm_table[1719] = 12'b000100_110000;
		logarithm_table[1720] = 12'b000100_110000;
		logarithm_table[1721] = 12'b000100_110000;
		logarithm_table[1722] = 12'b000100_110000;
		logarithm_table[1723] = 12'b000100_110000;
		logarithm_table[1724] = 12'b000100_110000;
		logarithm_table[1725] = 12'b000100_110000;
		logarithm_table[1726] = 12'b000100_110000;
		logarithm_table[1727] = 12'b000100_110000;
		logarithm_table[1728] = 12'b000100_110000;
		logarithm_table[1729] = 12'b000100_110000;
		logarithm_table[1730] = 12'b000100_110000;
		logarithm_table[1731] = 12'b000100_110000;
		logarithm_table[1732] = 12'b000100_110001;
		logarithm_table[1733] = 12'b000100_110001;
		logarithm_table[1734] = 12'b000100_110001;
		logarithm_table[1735] = 12'b000100_110001;
		logarithm_table[1736] = 12'b000100_110001;
		logarithm_table[1737] = 12'b000100_110001;
		logarithm_table[1738] = 12'b000100_110001;
		logarithm_table[1739] = 12'b000100_110001;
		logarithm_table[1740] = 12'b000100_110001;
		logarithm_table[1741] = 12'b000100_110001;
		logarithm_table[1742] = 12'b000100_110001;
		logarithm_table[1743] = 12'b000100_110001;
		logarithm_table[1744] = 12'b000100_110001;
		logarithm_table[1745] = 12'b000100_110001;
		logarithm_table[1746] = 12'b000100_110001;
		logarithm_table[1747] = 12'b000100_110001;
		logarithm_table[1748] = 12'b000100_110001;
		logarithm_table[1749] = 12'b000100_110001;
		logarithm_table[1750] = 12'b000100_110001;
		logarithm_table[1751] = 12'b000100_110010;
		logarithm_table[1752] = 12'b000100_110010;
		logarithm_table[1753] = 12'b000100_110010;
		logarithm_table[1754] = 12'b000100_110010;
		logarithm_table[1755] = 12'b000100_110010;
		logarithm_table[1756] = 12'b000100_110010;
		logarithm_table[1757] = 12'b000100_110010;
		logarithm_table[1758] = 12'b000100_110010;
		logarithm_table[1759] = 12'b000100_110010;
		logarithm_table[1760] = 12'b000100_110010;
		logarithm_table[1761] = 12'b000100_110010;
		logarithm_table[1762] = 12'b000100_110010;
		logarithm_table[1763] = 12'b000100_110010;
		logarithm_table[1764] = 12'b000100_110010;
		logarithm_table[1765] = 12'b000100_110010;
		logarithm_table[1766] = 12'b000100_110010;
		logarithm_table[1767] = 12'b000100_110010;
		logarithm_table[1768] = 12'b000100_110010;
		logarithm_table[1769] = 12'b000100_110010;
		logarithm_table[1770] = 12'b000100_110011;
		logarithm_table[1771] = 12'b000100_110011;
		logarithm_table[1772] = 12'b000100_110011;
		logarithm_table[1773] = 12'b000100_110011;
		logarithm_table[1774] = 12'b000100_110011;
		logarithm_table[1775] = 12'b000100_110011;
		logarithm_table[1776] = 12'b000100_110011;
		logarithm_table[1777] = 12'b000100_110011;
		logarithm_table[1778] = 12'b000100_110011;
		logarithm_table[1779] = 12'b000100_110011;
		logarithm_table[1780] = 12'b000100_110011;
		logarithm_table[1781] = 12'b000100_110011;
		logarithm_table[1782] = 12'b000100_110011;
		logarithm_table[1783] = 12'b000100_110011;
		logarithm_table[1784] = 12'b000100_110011;
		logarithm_table[1785] = 12'b000100_110011;
		logarithm_table[1786] = 12'b000100_110011;
		logarithm_table[1787] = 12'b000100_110011;
		logarithm_table[1788] = 12'b000100_110011;
		logarithm_table[1789] = 12'b000100_110100;
		logarithm_table[1790] = 12'b000100_110100;
		logarithm_table[1791] = 12'b000100_110100;
		logarithm_table[1792] = 12'b000100_110100;
		logarithm_table[1793] = 12'b000100_110100;
		logarithm_table[1794] = 12'b000100_110100;
		logarithm_table[1795] = 12'b000100_110100;
		logarithm_table[1796] = 12'b000100_110100;
		logarithm_table[1797] = 12'b000100_110100;
		logarithm_table[1798] = 12'b000100_110100;
		logarithm_table[1799] = 12'b000100_110100;
		logarithm_table[1800] = 12'b000100_110100;
		logarithm_table[1801] = 12'b000100_110100;
		logarithm_table[1802] = 12'b000100_110100;
		logarithm_table[1803] = 12'b000100_110100;
		logarithm_table[1804] = 12'b000100_110100;
		logarithm_table[1805] = 12'b000100_110100;
		logarithm_table[1806] = 12'b000100_110100;
		logarithm_table[1807] = 12'b000100_110100;
		logarithm_table[1808] = 12'b000100_110100;
		logarithm_table[1809] = 12'b000100_110101;
		logarithm_table[1810] = 12'b000100_110101;
		logarithm_table[1811] = 12'b000100_110101;
		logarithm_table[1812] = 12'b000100_110101;
		logarithm_table[1813] = 12'b000100_110101;
		logarithm_table[1814] = 12'b000100_110101;
		logarithm_table[1815] = 12'b000100_110101;
		logarithm_table[1816] = 12'b000100_110101;
		logarithm_table[1817] = 12'b000100_110101;
		logarithm_table[1818] = 12'b000100_110101;
		logarithm_table[1819] = 12'b000100_110101;
		logarithm_table[1820] = 12'b000100_110101;
		logarithm_table[1821] = 12'b000100_110101;
		logarithm_table[1822] = 12'b000100_110101;
		logarithm_table[1823] = 12'b000100_110101;
		logarithm_table[1824] = 12'b000100_110101;
		logarithm_table[1825] = 12'b000100_110101;
		logarithm_table[1826] = 12'b000100_110101;
		logarithm_table[1827] = 12'b000100_110101;
		logarithm_table[1828] = 12'b000100_110110;
		logarithm_table[1829] = 12'b000100_110110;
		logarithm_table[1830] = 12'b000100_110110;
		logarithm_table[1831] = 12'b000100_110110;
		logarithm_table[1832] = 12'b000100_110110;
		logarithm_table[1833] = 12'b000100_110110;
		logarithm_table[1834] = 12'b000100_110110;
		logarithm_table[1835] = 12'b000100_110110;
		logarithm_table[1836] = 12'b000100_110110;
		logarithm_table[1837] = 12'b000100_110110;
		logarithm_table[1838] = 12'b000100_110110;
		logarithm_table[1839] = 12'b000100_110110;
		logarithm_table[1840] = 12'b000100_110110;
		logarithm_table[1841] = 12'b000100_110110;
		logarithm_table[1842] = 12'b000100_110110;
		logarithm_table[1843] = 12'b000100_110110;
		logarithm_table[1844] = 12'b000100_110110;
		logarithm_table[1845] = 12'b000100_110110;
		logarithm_table[1846] = 12'b000100_110110;
		logarithm_table[1847] = 12'b000100_110110;
		logarithm_table[1848] = 12'b000100_110111;
		logarithm_table[1849] = 12'b000100_110111;
		logarithm_table[1850] = 12'b000100_110111;
		logarithm_table[1851] = 12'b000100_110111;
		logarithm_table[1852] = 12'b000100_110111;
		logarithm_table[1853] = 12'b000100_110111;
		logarithm_table[1854] = 12'b000100_110111;
		logarithm_table[1855] = 12'b000100_110111;
		logarithm_table[1856] = 12'b000100_110111;
		logarithm_table[1857] = 12'b000100_110111;
		logarithm_table[1858] = 12'b000100_110111;
		logarithm_table[1859] = 12'b000100_110111;
		logarithm_table[1860] = 12'b000100_110111;
		logarithm_table[1861] = 12'b000100_110111;
		logarithm_table[1862] = 12'b000100_110111;
		logarithm_table[1863] = 12'b000100_110111;
		logarithm_table[1864] = 12'b000100_110111;
		logarithm_table[1865] = 12'b000100_110111;
		logarithm_table[1866] = 12'b000100_110111;
		logarithm_table[1867] = 12'b000100_110111;
		logarithm_table[1868] = 12'b000100_111000;
		logarithm_table[1869] = 12'b000100_111000;
		logarithm_table[1870] = 12'b000100_111000;
		logarithm_table[1871] = 12'b000100_111000;
		logarithm_table[1872] = 12'b000100_111000;
		logarithm_table[1873] = 12'b000100_111000;
		logarithm_table[1874] = 12'b000100_111000;
		logarithm_table[1875] = 12'b000100_111000;
		logarithm_table[1876] = 12'b000100_111000;
		logarithm_table[1877] = 12'b000100_111000;
		logarithm_table[1878] = 12'b000100_111000;
		logarithm_table[1879] = 12'b000100_111000;
		logarithm_table[1880] = 12'b000100_111000;
		logarithm_table[1881] = 12'b000100_111000;
		logarithm_table[1882] = 12'b000100_111000;
		logarithm_table[1883] = 12'b000100_111000;
		logarithm_table[1884] = 12'b000100_111000;
		logarithm_table[1885] = 12'b000100_111000;
		logarithm_table[1886] = 12'b000100_111000;
		logarithm_table[1887] = 12'b000100_111000;
		logarithm_table[1888] = 12'b000100_111000;
		logarithm_table[1889] = 12'b000100_111001;
		logarithm_table[1890] = 12'b000100_111001;
		logarithm_table[1891] = 12'b000100_111001;
		logarithm_table[1892] = 12'b000100_111001;
		logarithm_table[1893] = 12'b000100_111001;
		logarithm_table[1894] = 12'b000100_111001;
		logarithm_table[1895] = 12'b000100_111001;
		logarithm_table[1896] = 12'b000100_111001;
		logarithm_table[1897] = 12'b000100_111001;
		logarithm_table[1898] = 12'b000100_111001;
		logarithm_table[1899] = 12'b000100_111001;
		logarithm_table[1900] = 12'b000100_111001;
		logarithm_table[1901] = 12'b000100_111001;
		logarithm_table[1902] = 12'b000100_111001;
		logarithm_table[1903] = 12'b000100_111001;
		logarithm_table[1904] = 12'b000100_111001;
		logarithm_table[1905] = 12'b000100_111001;
		logarithm_table[1906] = 12'b000100_111001;
		logarithm_table[1907] = 12'b000100_111001;
		logarithm_table[1908] = 12'b000100_111001;
		logarithm_table[1909] = 12'b000100_111010;
		logarithm_table[1910] = 12'b000100_111010;
		logarithm_table[1911] = 12'b000100_111010;
		logarithm_table[1912] = 12'b000100_111010;
		logarithm_table[1913] = 12'b000100_111010;
		logarithm_table[1914] = 12'b000100_111010;
		logarithm_table[1915] = 12'b000100_111010;
		logarithm_table[1916] = 12'b000100_111010;
		logarithm_table[1917] = 12'b000100_111010;
		logarithm_table[1918] = 12'b000100_111010;
		logarithm_table[1919] = 12'b000100_111010;
		logarithm_table[1920] = 12'b000100_111010;
		logarithm_table[1921] = 12'b000100_111010;
		logarithm_table[1922] = 12'b000100_111010;
		logarithm_table[1923] = 12'b000100_111010;
		logarithm_table[1924] = 12'b000100_111010;
		logarithm_table[1925] = 12'b000100_111010;
		logarithm_table[1926] = 12'b000100_111010;
		logarithm_table[1927] = 12'b000100_111010;
		logarithm_table[1928] = 12'b000100_111010;
		logarithm_table[1929] = 12'b000100_111010;
		logarithm_table[1930] = 12'b000100_111011;
		logarithm_table[1931] = 12'b000100_111011;
		logarithm_table[1932] = 12'b000100_111011;
		logarithm_table[1933] = 12'b000100_111011;
		logarithm_table[1934] = 12'b000100_111011;
		logarithm_table[1935] = 12'b000100_111011;
		logarithm_table[1936] = 12'b000100_111011;
		logarithm_table[1937] = 12'b000100_111011;
		logarithm_table[1938] = 12'b000100_111011;
		logarithm_table[1939] = 12'b000100_111011;
		logarithm_table[1940] = 12'b000100_111011;
		logarithm_table[1941] = 12'b000100_111011;
		logarithm_table[1942] = 12'b000100_111011;
		logarithm_table[1943] = 12'b000100_111011;
		logarithm_table[1944] = 12'b000100_111011;
		logarithm_table[1945] = 12'b000100_111011;
		logarithm_table[1946] = 12'b000100_111011;
		logarithm_table[1947] = 12'b000100_111011;
		logarithm_table[1948] = 12'b000100_111011;
		logarithm_table[1949] = 12'b000100_111011;
		logarithm_table[1950] = 12'b000100_111011;
		logarithm_table[1951] = 12'b000100_111100;
		logarithm_table[1952] = 12'b000100_111100;
		logarithm_table[1953] = 12'b000100_111100;
		logarithm_table[1954] = 12'b000100_111100;
		logarithm_table[1955] = 12'b000100_111100;
		logarithm_table[1956] = 12'b000100_111100;
		logarithm_table[1957] = 12'b000100_111100;
		logarithm_table[1958] = 12'b000100_111100;
		logarithm_table[1959] = 12'b000100_111100;
		logarithm_table[1960] = 12'b000100_111100;
		logarithm_table[1961] = 12'b000100_111100;
		logarithm_table[1962] = 12'b000100_111100;
		logarithm_table[1963] = 12'b000100_111100;
		logarithm_table[1964] = 12'b000100_111100;
		logarithm_table[1965] = 12'b000100_111100;
		logarithm_table[1966] = 12'b000100_111100;
		logarithm_table[1967] = 12'b000100_111100;
		logarithm_table[1968] = 12'b000100_111100;
		logarithm_table[1969] = 12'b000100_111100;
		logarithm_table[1970] = 12'b000100_111100;
		logarithm_table[1971] = 12'b000100_111100;
		logarithm_table[1972] = 12'b000100_111101;
		logarithm_table[1973] = 12'b000100_111101;
		logarithm_table[1974] = 12'b000100_111101;
		logarithm_table[1975] = 12'b000100_111101;
		logarithm_table[1976] = 12'b000100_111101;
		logarithm_table[1977] = 12'b000100_111101;
		logarithm_table[1978] = 12'b000100_111101;
		logarithm_table[1979] = 12'b000100_111101;
		logarithm_table[1980] = 12'b000100_111101;
		logarithm_table[1981] = 12'b000100_111101;
		logarithm_table[1982] = 12'b000100_111101;
		logarithm_table[1983] = 12'b000100_111101;
		logarithm_table[1984] = 12'b000100_111101;
		logarithm_table[1985] = 12'b000100_111101;
		logarithm_table[1986] = 12'b000100_111101;
		logarithm_table[1987] = 12'b000100_111101;
		logarithm_table[1988] = 12'b000100_111101;
		logarithm_table[1989] = 12'b000100_111101;
		logarithm_table[1990] = 12'b000100_111101;
		logarithm_table[1991] = 12'b000100_111101;
		logarithm_table[1992] = 12'b000100_111101;
		logarithm_table[1993] = 12'b000100_111101;
		logarithm_table[1994] = 12'b000100_111110;
		logarithm_table[1995] = 12'b000100_111110;
		logarithm_table[1996] = 12'b000100_111110;
		logarithm_table[1997] = 12'b000100_111110;
		logarithm_table[1998] = 12'b000100_111110;
		logarithm_table[1999] = 12'b000100_111110;
		logarithm_table[2000] = 12'b000100_111110;
		logarithm_table[2001] = 12'b000100_111110;
		logarithm_table[2002] = 12'b000100_111110;
		logarithm_table[2003] = 12'b000100_111110;
		logarithm_table[2004] = 12'b000100_111110;
		logarithm_table[2005] = 12'b000100_111110;
		logarithm_table[2006] = 12'b000100_111110;
		logarithm_table[2007] = 12'b000100_111110;
		logarithm_table[2008] = 12'b000100_111110;
		logarithm_table[2009] = 12'b000100_111110;
		logarithm_table[2010] = 12'b000100_111110;
		logarithm_table[2011] = 12'b000100_111110;
		logarithm_table[2012] = 12'b000100_111110;
		logarithm_table[2013] = 12'b000100_111110;
		logarithm_table[2014] = 12'b000100_111110;
		logarithm_table[2015] = 12'b000100_111111;
		logarithm_table[2016] = 12'b000100_111111;
		logarithm_table[2017] = 12'b000100_111111;
		logarithm_table[2018] = 12'b000100_111111;
		logarithm_table[2019] = 12'b000100_111111;
		logarithm_table[2020] = 12'b000100_111111;
		logarithm_table[2021] = 12'b000100_111111;
		logarithm_table[2022] = 12'b000100_111111;
		logarithm_table[2023] = 12'b000100_111111;
		logarithm_table[2024] = 12'b000100_111111;
		logarithm_table[2025] = 12'b000100_111111;
		logarithm_table[2026] = 12'b000100_111111;
		logarithm_table[2027] = 12'b000100_111111;
		logarithm_table[2028] = 12'b000100_111111;
		logarithm_table[2029] = 12'b000100_111111;
		logarithm_table[2030] = 12'b000100_111111;
		logarithm_table[2031] = 12'b000100_111111;
		logarithm_table[2032] = 12'b000100_111111;
		logarithm_table[2033] = 12'b000100_111111;
		logarithm_table[2034] = 12'b000100_111111;
		logarithm_table[2035] = 12'b000100_111111;
		logarithm_table[2036] = 12'b000100_111111;
		logarithm_table[2037] = 12'b000101_000000;
		logarithm_table[2038] = 12'b000101_000000;
		logarithm_table[2039] = 12'b000101_000000;
		logarithm_table[2040] = 12'b000101_000000;
		logarithm_table[2041] = 12'b000101_000000;
		logarithm_table[2042] = 12'b000101_000000;
		logarithm_table[2043] = 12'b000101_000000;
		logarithm_table[2044] = 12'b000101_000000;
		logarithm_table[2045] = 12'b000101_000000;
		logarithm_table[2046] = 12'b000101_000000;
		logarithm_table[2047] = 12'b000101_000000;
		Dminus[1] = 12'b111110_100001;
		Dminus[2] = 12'b111110_100010;
		Dminus[3] = 12'b111110_100011;
		Dminus[4] = 12'b111110_100100;
		Dminus[5] = 12'b111110_100101;
		Dminus[6] = 12'b111110_100110;
		Dminus[7] = 12'b111110_100111;
		Dminus[8] = 12'b111110_101000;
		Dminus[9] = 12'b111110_101001;
		Dminus[10] = 12'b111110_101010;
		Dminus[11] = 12'b111110_101011;
		Dminus[12] = 12'b111110_101100;
		Dminus[13] = 12'b111110_101101;
		Dminus[14] = 12'b111110_101110;
		Dminus[15] = 12'b111110_101110;
		Dminus[16] = 12'b111110_101111;
		Dminus[17] = 12'b111110_110000;
		Dminus[18] = 12'b111110_110001;
		Dminus[19] = 12'b111110_110010;
		Dminus[20] = 12'b111110_110011;
		Dminus[21] = 12'b111110_110100;
		Dminus[22] = 12'b111110_110100;
		Dminus[23] = 12'b111110_110101;
		Dminus[24] = 12'b111110_110110;
		Dminus[25] = 12'b111110_110111;
		Dminus[26] = 12'b111110_111000;
		Dminus[27] = 12'b111110_111000;
		Dminus[28] = 12'b111110_111001;
		Dminus[29] = 12'b111110_111010;
		Dminus[30] = 12'b111110_111011;
		Dminus[31] = 12'b111110_111011;
		Dminus[32] = 12'b111110_111100;
		Dminus[33] = 12'b111110_111101;
		Dminus[34] = 12'b111110_111110;
		Dminus[35] = 12'b111110_111110;
		Dminus[36] = 12'b111110_111111;
		Dminus[37] = 12'b111111_000000;
		Dminus[38] = 12'b111111_000000;
		Dminus[39] = 12'b111111_000001;
		Dminus[40] = 12'b111111_000010;
		Dminus[41] = 12'b111111_000010;
		Dminus[42] = 12'b111111_000011;
		Dminus[43] = 12'b111111_000100;
		Dminus[44] = 12'b111111_000100;
		Dminus[45] = 12'b111111_000101;
		Dminus[46] = 12'b111111_000110;
		Dminus[47] = 12'b111111_000110;
		Dminus[48] = 12'b111111_000111;
		Dminus[49] = 12'b111111_001000;
		Dminus[50] = 12'b111111_001000;
		Dminus[51] = 12'b111111_001001;
		Dminus[52] = 12'b111111_001001;
		Dminus[53] = 12'b111111_001010;
		Dminus[54] = 12'b111111_001011;
		Dminus[55] = 12'b111111_001011;
		Dminus[56] = 12'b111111_001100;
		Dminus[57] = 12'b111111_001100;
		Dminus[58] = 12'b111111_001101;
		Dminus[59] = 12'b111111_001101;
		Dminus[60] = 12'b111111_001110;
		Dminus[61] = 12'b111111_001110;
		Dminus[62] = 12'b111111_001111;
		Dminus[63] = 12'b111111_001111;
		Dminus[64] = 12'b111111_010000;
		Dminus[65] = 12'b111111_010001;
		Dminus[66] = 12'b111111_010001;
		Dminus[67] = 12'b111111_010010;
		Dminus[68] = 12'b111111_010010;
		Dminus[69] = 12'b111111_010011;
		Dminus[70] = 12'b111111_010011;
		Dminus[71] = 12'b111111_010100;
		Dminus[72] = 12'b111111_010100;
		Dminus[73] = 12'b111111_010100;
		Dminus[74] = 12'b111111_010101;
		Dminus[75] = 12'b111111_010101;
		Dminus[76] = 12'b111111_010110;
		Dminus[77] = 12'b111111_010110;
		Dminus[78] = 12'b111111_010111;
		Dminus[79] = 12'b111111_010111;
		Dminus[80] = 12'b111111_011000;
		Dminus[81] = 12'b111111_011000;
		Dminus[82] = 12'b111111_011001;
		Dminus[83] = 12'b111111_011001;
		Dminus[84] = 12'b111111_011001;
		Dminus[85] = 12'b111111_011010;
		Dminus[86] = 12'b111111_011010;
		Dminus[87] = 12'b111111_011011;
		Dminus[88] = 12'b111111_011011;
		Dminus[89] = 12'b111111_011011;
		Dminus[90] = 12'b111111_011100;
		Dminus[91] = 12'b111111_011100;
		Dminus[92] = 12'b111111_011101;
		Dminus[93] = 12'b111111_011101;
		Dminus[94] = 12'b111111_011101;
		Dminus[95] = 12'b111111_011110;
		Dminus[96] = 12'b111111_011110;
		Dminus[97] = 12'b111111_011110;
		Dminus[98] = 12'b111111_011111;
		Dminus[99] = 12'b111111_011111;
		Dminus[100] = 12'b111111_011111;
		Dminus[101] = 12'b111111_100000;
		Dminus[102] = 12'b111111_100000;
		Dminus[103] = 12'b111111_100001;
		Dminus[104] = 12'b111111_100001;
		Dminus[105] = 12'b111111_100001;
		Dminus[106] = 12'b111111_100010;
		Dminus[107] = 12'b111111_100010;
		Dminus[108] = 12'b111111_100010;
		Dminus[109] = 12'b111111_100011;
		Dminus[110] = 12'b111111_100011;
		Dminus[111] = 12'b111111_100011;
		Dminus[112] = 12'b111111_100011;
		Dminus[113] = 12'b111111_100100;
		Dminus[114] = 12'b111111_100100;
		Dminus[115] = 12'b111111_100100;
		Dminus[116] = 12'b111111_100101;
		Dminus[117] = 12'b111111_100101;
		Dminus[118] = 12'b111111_100101;
		Dminus[119] = 12'b111111_100110;
		Dminus[120] = 12'b111111_100110;
		Dminus[121] = 12'b111111_100110;
		Dminus[122] = 12'b111111_100110;
		Dminus[123] = 12'b111111_100111;
		Dminus[124] = 12'b111111_100111;
		Dminus[125] = 12'b111111_100111;
		Dminus[126] = 12'b111111_100111;
		Dminus[127] = 12'b111111_101000;
		Dminus[128] = 12'b111111_101000;
		Dminus[129] = 12'b111111_101000;
		Dminus[130] = 12'b111111_101001;
		Dminus[131] = 12'b111111_101001;
		Dminus[132] = 12'b111111_101001;
		Dminus[133] = 12'b111111_101001;
		Dminus[134] = 12'b111111_101010;
		Dminus[135] = 12'b111111_101010;
		Dminus[136] = 12'b111111_101010;
		Dminus[137] = 12'b111111_101010;
		Dminus[138] = 12'b111111_101010;
		Dminus[139] = 12'b111111_101011;
		Dminus[140] = 12'b111111_101011;
		Dminus[141] = 12'b111111_101011;
		Dminus[142] = 12'b111111_101011;
		Dminus[143] = 12'b111111_101100;
		Dminus[144] = 12'b111111_101100;
		Dminus[145] = 12'b111111_101100;
		Dminus[146] = 12'b111111_101100;
		Dminus[147] = 12'b111111_101100;
		Dminus[148] = 12'b111111_101101;
		Dminus[149] = 12'b111111_101101;
		Dminus[150] = 12'b111111_101101;
		Dminus[151] = 12'b111111_101101;
		Dminus[152] = 12'b111111_101101;
		Dminus[153] = 12'b111111_101110;
		Dminus[154] = 12'b111111_101110;
		Dminus[155] = 12'b111111_101110;
		Dminus[156] = 12'b111111_101110;
		Dminus[157] = 12'b111111_101110;
		Dminus[158] = 12'b111111_101111;
		Dminus[159] = 12'b111111_101111;
		Dminus[160] = 12'b111111_101111;
		Dminus[161] = 12'b111111_101111;
		Dminus[162] = 12'b111111_101111;
		Dminus[163] = 12'b111111_110000;
		Dminus[164] = 12'b111111_110000;
		Dminus[165] = 12'b111111_110000;
		Dminus[166] = 12'b111111_110000;
		Dminus[167] = 12'b111111_110000;
		Dminus[168] = 12'b111111_110000;
		Dminus[169] = 12'b111111_110001;
		Dminus[170] = 12'b111111_110001;
		Dminus[171] = 12'b111111_110001;
		Dminus[172] = 12'b111111_110001;
		Dminus[173] = 12'b111111_110001;
		Dminus[174] = 12'b111111_110001;
		Dminus[175] = 12'b111111_110010;
		Dminus[176] = 12'b111111_110010;
		Dminus[177] = 12'b111111_110010;
		Dminus[178] = 12'b111111_110010;
		Dminus[179] = 12'b111111_110010;
		Dminus[180] = 12'b111111_110010;
		Dminus[181] = 12'b111111_110010;
		Dminus[182] = 12'b111111_110011;
		Dminus[183] = 12'b111111_110011;
		Dminus[184] = 12'b111111_110011;
		Dminus[185] = 12'b111111_110011;
		Dminus[186] = 12'b111111_110011;
		Dminus[187] = 12'b111111_110011;
		Dminus[188] = 12'b111111_110011;
		Dminus[189] = 12'b111111_110100;
		Dminus[190] = 12'b111111_110100;
		Dminus[191] = 12'b111111_110100;
		Dminus[192] = 12'b111111_110100;
		Dminus[193] = 12'b111111_110100;
		Dminus[194] = 12'b111111_110100;
		Dminus[195] = 12'b111111_110100;
		Dminus[196] = 12'b111111_110101;
		Dminus[197] = 12'b111111_110101;
		Dminus[198] = 12'b111111_110101;
		Dminus[199] = 12'b111111_110101;
		Dminus[200] = 12'b111111_110101;
		Dminus[201] = 12'b111111_110101;
		Dminus[202] = 12'b111111_110101;
		Dminus[203] = 12'b111111_110101;
		Dminus[204] = 12'b111111_110101;
		Dminus[205] = 12'b111111_110110;
		Dminus[206] = 12'b111111_110110;
		Dminus[207] = 12'b111111_110110;
		Dminus[208] = 12'b111111_110110;
		Dminus[209] = 12'b111111_110110;
		Dminus[210] = 12'b111111_110110;
		Dminus[211] = 12'b111111_110110;
		Dminus[212] = 12'b111111_110110;
		Dminus[213] = 12'b111111_110110;
		Dminus[214] = 12'b111111_110111;
		Dminus[215] = 12'b111111_110111;
		Dminus[216] = 12'b111111_110111;
		Dminus[217] = 12'b111111_110111;
		Dminus[218] = 12'b111111_110111;
		Dminus[219] = 12'b111111_110111;
		Dminus[220] = 12'b111111_110111;
		Dminus[221] = 12'b111111_110111;
		Dminus[222] = 12'b111111_110111;
		Dminus[223] = 12'b111111_110111;
		Dminus[224] = 12'b111111_111000;
		Dminus[225] = 12'b111111_111000;
		Dminus[226] = 12'b111111_111000;
		Dminus[227] = 12'b111111_111000;
		Dminus[228] = 12'b111111_111000;
		Dminus[229] = 12'b111111_111000;
		Dminus[230] = 12'b111111_111000;
		Dminus[231] = 12'b111111_111000;
		Dminus[232] = 12'b111111_111000;
		Dminus[233] = 12'b111111_111000;
		Dminus[234] = 12'b111111_111000;
		Dminus[235] = 12'b111111_111000;
		Dminus[236] = 12'b111111_111001;
		Dminus[237] = 12'b111111_111001;
		Dminus[238] = 12'b111111_111001;
		Dminus[239] = 12'b111111_111001;
		Dminus[240] = 12'b111111_111001;
		Dminus[241] = 12'b111111_111001;
		Dminus[242] = 12'b111111_111001;
		Dminus[243] = 12'b111111_111001;
		Dminus[244] = 12'b111111_111001;
		Dminus[245] = 12'b111111_111001;
		Dminus[246] = 12'b111111_111001;
		Dminus[247] = 12'b111111_111001;
		Dminus[248] = 12'b111111_111001;
		Dminus[249] = 12'b111111_111010;
		Dminus[250] = 12'b111111_111010;
		Dminus[251] = 12'b111111_111010;
		Dminus[252] = 12'b111111_111010;
		Dminus[253] = 12'b111111_111010;
		Dminus[254] = 12'b111111_111010;
		Dminus[255] = 12'b111111_111010;
		Dminus[256] = 12'b111111_111010;
		Dminus[257] = 12'b111111_111010;
		Dminus[258] = 12'b111111_111010;
		Dminus[259] = 12'b111111_111010;
		Dminus[260] = 12'b111111_111010;
		Dminus[261] = 12'b111111_111010;
		Dminus[262] = 12'b111111_111010;
		Dminus[263] = 12'b111111_111010;
		Dminus[264] = 12'b111111_111010;
		Dminus[265] = 12'b111111_111011;
		Dminus[266] = 12'b111111_111011;
		Dminus[267] = 12'b111111_111011;
		Dminus[268] = 12'b111111_111011;
		Dminus[269] = 12'b111111_111011;
		Dminus[270] = 12'b111111_111011;
		Dminus[271] = 12'b111111_111011;
		Dminus[272] = 12'b111111_111011;
		Dminus[273] = 12'b111111_111011;
		Dminus[274] = 12'b111111_111011;
		Dminus[275] = 12'b111111_111011;
		Dminus[276] = 12'b111111_111011;
		Dminus[277] = 12'b111111_111011;
		Dminus[278] = 12'b111111_111011;
		Dminus[279] = 12'b111111_111011;
		Dminus[280] = 12'b111111_111011;
		Dminus[281] = 12'b111111_111011;
		Dminus[282] = 12'b111111_111011;
		Dminus[283] = 12'b111111_111100;
		Dminus[284] = 12'b111111_111100;
		Dminus[285] = 12'b111111_111100;
		Dminus[286] = 12'b111111_111100;
		Dminus[287] = 12'b111111_111100;
		Dminus[288] = 12'b111111_111100;
		Dminus[289] = 12'b111111_111100;
		Dminus[290] = 12'b111111_111100;
		Dminus[291] = 12'b111111_111100;
		Dminus[292] = 12'b111111_111100;
		Dminus[293] = 12'b111111_111100;
		Dminus[294] = 12'b111111_111100;
		Dminus[295] = 12'b111111_111100;
		Dminus[296] = 12'b111111_111100;
		Dminus[297] = 12'b111111_111100;
		Dminus[298] = 12'b111111_111100;
		Dminus[299] = 12'b111111_111100;
		Dminus[300] = 12'b111111_111100;
		Dminus[301] = 12'b111111_111100;
		Dminus[302] = 12'b111111_111100;
		Dminus[303] = 12'b111111_111100;
		Dminus[304] = 12'b111111_111100;
		Dminus[305] = 12'b111111_111100;
		Dminus[306] = 12'b111111_111101;
		Dminus[307] = 12'b111111_111101;
		Dminus[308] = 12'b111111_111101;
		Dminus[309] = 12'b111111_111101;
		Dminus[310] = 12'b111111_111101;
		Dminus[311] = 12'b111111_111101;
		Dminus[312] = 12'b111111_111101;
		Dminus[313] = 12'b111111_111101;
		Dminus[314] = 12'b111111_111101;
		Dminus[315] = 12'b111111_111101;
		Dminus[316] = 12'b111111_111101;
		Dminus[317] = 12'b111111_111101;
		Dminus[318] = 12'b111111_111101;
		Dminus[319] = 12'b111111_111101;
		Dminus[320] = 12'b111111_111101;
		Dminus[321] = 12'b111111_111101;
		Dminus[322] = 12'b111111_111101;
		Dminus[323] = 12'b111111_111101;
		Dminus[324] = 12'b111111_111101;
		Dminus[325] = 12'b111111_111101;
		Dminus[326] = 12'b111111_111101;
		Dminus[327] = 12'b111111_111101;
		Dminus[328] = 12'b111111_111101;
		Dminus[329] = 12'b111111_111101;
		Dminus[330] = 12'b111111_111101;
		Dminus[331] = 12'b111111_111101;
		Dminus[332] = 12'b111111_111101;
		Dminus[333] = 12'b111111_111101;
		Dminus[334] = 12'b111111_111101;
		Dminus[335] = 12'b111111_111101;
		Dminus[336] = 12'b111111_111101;
		Dminus[337] = 12'b111111_111110;
		Dminus[338] = 12'b111111_111110;
		Dminus[339] = 12'b111111_111110;
		Dminus[340] = 12'b111111_111110;
		Dminus[341] = 12'b111111_111110;
		Dminus[342] = 12'b111111_111110;
		Dminus[343] = 12'b111111_111110;
		Dminus[344] = 12'b111111_111110;
		Dminus[345] = 12'b111111_111110;
		Dminus[346] = 12'b111111_111110;
		Dminus[347] = 12'b111111_111110;
		Dminus[348] = 12'b111111_111110;
		Dminus[349] = 12'b111111_111110;
		Dminus[350] = 12'b111111_111110;
		Dminus[351] = 12'b111111_111110;
		Dminus[352] = 12'b111111_111110;
		Dminus[353] = 12'b111111_111110;
		Dminus[354] = 12'b111111_111110;
		Dminus[355] = 12'b111111_111110;
		Dminus[356] = 12'b111111_111110;
		Dminus[357] = 12'b111111_111110;
		Dminus[358] = 12'b111111_111110;
		Dminus[359] = 12'b111111_111110;
		Dminus[360] = 12'b111111_111110;
		Dminus[361] = 12'b111111_111110;
		Dminus[362] = 12'b111111_111110;
		Dminus[363] = 12'b111111_111110;
		Dminus[364] = 12'b111111_111110;
		Dminus[365] = 12'b111111_111110;
		Dminus[366] = 12'b111111_111110;
		Dminus[367] = 12'b111111_111110;
		Dminus[368] = 12'b111111_111110;
		Dminus[369] = 12'b111111_111110;
		Dminus[370] = 12'b111111_111110;
		Dminus[371] = 12'b111111_111110;
		Dminus[372] = 12'b111111_111110;
		Dminus[373] = 12'b111111_111110;
		Dminus[374] = 12'b111111_111110;
		Dminus[375] = 12'b111111_111110;
		Dminus[376] = 12'b111111_111110;
		Dminus[377] = 12'b111111_111110;
		Dminus[378] = 12'b111111_111110;
		Dminus[379] = 12'b111111_111110;
		Dminus[380] = 12'b111111_111110;
		Dminus[381] = 12'b111111_111110;
		Dminus[382] = 12'b111111_111110;
		Dminus[383] = 12'b111111_111110;
		Dminus[384] = 12'b111111_111110;
		Dminus[385] = 12'b111111_111111;
		Dminus[386] = 12'b111111_111111;
		Dminus[387] = 12'b111111_111111;
		Dminus[388] = 12'b111111_111111;
		Dminus[389] = 12'b111111_111111;
		Dminus[390] = 12'b111111_111111;
		Dminus[391] = 12'b111111_111111;
		Dminus[392] = 12'b111111_111111;
		Dminus[393] = 12'b111111_111111;
		Dminus[394] = 12'b111111_111111;
		Dminus[395] = 12'b111111_111111;
		Dminus[396] = 12'b111111_111111;
		Dminus[397] = 12'b111111_111111;
		Dminus[398] = 12'b111111_111111;
		Dminus[399] = 12'b111111_111111;
		Dminus[400] = 12'b111111_111111;
		Dminus[401] = 12'b111111_111111;
		Dminus[402] = 12'b111111_111111;
		Dminus[403] = 12'b111111_111111;
		Dminus[404] = 12'b111111_111111;
		Dminus[405] = 12'b111111_111111;
		Dminus[406] = 12'b111111_111111;
		Dminus[407] = 12'b111111_111111;
		Dminus[408] = 12'b111111_111111;
		Dminus[409] = 12'b111111_111111;
		Dminus[410] = 12'b111111_111111;
		Dminus[411] = 12'b111111_111111;
		Dminus[412] = 12'b111111_111111;
		Dminus[413] = 12'b111111_111111;
		Dminus[414] = 12'b111111_111111;
		Dminus[415] = 12'b111111_111111;
		Dminus[416] = 12'b111111_111111;
		Dminus[417] = 12'b111111_111111;
		Dminus[418] = 12'b111111_111111;
		Dminus[419] = 12'b111111_111111;
		Dminus[420] = 12'b111111_111111;
		Dminus[421] = 12'b111111_111111;
		Dminus[422] = 12'b111111_111111;
		Dminus[423] = 12'b111111_111111;
		Dminus[424] = 12'b111111_111111;
		Dminus[425] = 12'b111111_111111;
		Dminus[426] = 12'b111111_111111;
		Dminus[427] = 12'b111111_111111;
		Dminus[428] = 12'b111111_111111;
		Dminus[429] = 12'b111111_111111;
		Dminus[430] = 12'b111111_111111;
		Dminus[431] = 12'b111111_111111;
		Dminus[432] = 12'b111111_111111;
		Dminus[433] = 12'b111111_111111;
		Dminus[434] = 12'b111111_111111;
		Dminus[435] = 12'b111111_111111;
		Dminus[436] = 12'b111111_111111;
		Dminus[437] = 12'b111111_111111;
		Dminus[438] = 12'b111111_111111;
		Dminus[439] = 12'b111111_111111;
		Dminus[440] = 12'b111111_111111;
		Dminus[441] = 12'b111111_111111;
		Dminus[442] = 12'b111111_111111;
		Dminus[443] = 12'b111111_111111;
		Dminus[444] = 12'b111111_111111;
		Dminus[445] = 12'b111111_111111;
		Dminus[446] = 12'b111111_111111;
		Dminus[447] = 12'b111111_111111;
		Dminus[448] = 12'b111111_111111;
		Dminus[449] = 12'b111111_111111;
		Dminus[450] = 12'b111111_111111;
		Dminus[451] = 12'b111111_111111;
		Dminus[452] = 12'b111111_111111;
		Dminus[453] = 12'b111111_111111;
		Dminus[454] = 12'b111111_111111;
		Dminus[455] = 12'b111111_111111;
		Dminus[456] = 12'b111111_111111;
		Dminus[457] = 12'b111111_111111;
		Dminus[458] = 12'b111111_111111;
		Dminus[459] = 12'b111111_111111;
		Dminus[460] = 12'b111111_111111;
		Dminus[461] = 12'b111111_111111;
		Dminus[462] = 12'b111111_111111;
		Dminus[463] = 12'b111111_111111;
		Dminus[464] = 12'b111111_111111;
		Dminus[465] = 12'b111111_111111;
		Dminus[466] = 12'b111111_111111;
		Dminus[467] = 12'b111111_111111;
		Dminus[468] = 12'b111111_111111;
		Dminus[469] = 12'b111111_111111;
		Dminus[470] = 12'b111111_111111;
		Dminus[471] = 12'b111111_111111;
		Dminus[472] = 12'b111111_111111;
		Dminus[473] = 12'b111111_111111;
		Dminus[474] = 12'b111111_111111;
		Dminus[475] = 12'b111111_111111;
		Dminus[476] = 12'b111111_111111;
		Dminus[477] = 12'b111111_111111;
		Dminus[478] = 12'b111111_111111;
		Dminus[479] = 12'b111111_111111;
		Dminus[480] = 12'b111111_111111;
		Dminus[481] = 12'b111111_111111;
		Dminus[482] = 12'b111111_111111;
		Dminus[483] = 12'b111111_111111;
		Dminus[484] = 12'b111111_111111;
		Dminus[485] = 12'b111111_111111;
		Dminus[486] = 12'b000000_000000;
		Dminus[487] = 12'b000000_000000;
		Dminus[488] = 12'b000000_000000;
		Dminus[489] = 12'b000000_000000;
		Dminus[490] = 12'b000000_000000;
		Dminus[491] = 12'b000000_000000;
		Dminus[492] = 12'b000000_000000;
		Dminus[493] = 12'b000000_000000;
		Dminus[494] = 12'b000000_000000;
		Dminus[495] = 12'b000000_000000;
		Dminus[496] = 12'b000000_000000;
		Dminus[497] = 12'b000000_000000;
		Dminus[498] = 12'b000000_000000;
		Dminus[499] = 12'b000000_000000;
		Dminus[500] = 12'b000000_000000;
		Dminus[501] = 12'b000000_000000;
		Dminus[502] = 12'b000000_000000;
		Dminus[503] = 12'b000000_000000;
		Dminus[504] = 12'b000000_000000;
		Dminus[505] = 12'b000000_000000;
		Dminus[506] = 12'b000000_000000;
		Dminus[507] = 12'b000000_000000;
		Dminus[508] = 12'b000000_000000;
		Dminus[509] = 12'b000000_000000;
		Dminus[510] = 12'b000000_000000;
		Dminus[511] = 12'b000000_000000;
		Dminus[512] = 12'b000000_000000;
		Dminus[513] = 12'b000000_000000;
		Dminus[514] = 12'b000000_000000;
		Dminus[515] = 12'b000000_000000;
		Dminus[516] = 12'b000000_000000;
		Dminus[517] = 12'b000000_000000;
		Dminus[518] = 12'b000000_000000;
		Dminus[519] = 12'b000000_000000;
		Dminus[520] = 12'b000000_000000;
		Dminus[521] = 12'b000000_000000;
		Dminus[522] = 12'b000000_000000;
		Dminus[523] = 12'b000000_000000;
		Dminus[524] = 12'b000000_000000;
		Dminus[525] = 12'b000000_000000;
		Dminus[526] = 12'b000000_000000;
		Dminus[527] = 12'b000000_000000;
		Dminus[528] = 12'b000000_000000;
		Dminus[529] = 12'b000000_000000;
		Dminus[530] = 12'b000000_000000;
		Dminus[531] = 12'b000000_000000;
		Dminus[532] = 12'b000000_000000;
		Dminus[533] = 12'b000000_000000;
		Dminus[534] = 12'b000000_000000;
		Dminus[535] = 12'b000000_000000;
		Dminus[536] = 12'b000000_000000;
		Dminus[537] = 12'b000000_000000;
		Dminus[538] = 12'b000000_000000;
		Dminus[539] = 12'b000000_000000;
		Dminus[540] = 12'b000000_000000;
		Dminus[541] = 12'b000000_000000;
		Dminus[542] = 12'b000000_000000;
		Dminus[543] = 12'b000000_000000;
		Dminus[544] = 12'b000000_000000;
		Dminus[545] = 12'b000000_000000;
		Dminus[546] = 12'b000000_000000;
		Dminus[547] = 12'b000000_000000;
		Dminus[548] = 12'b000000_000000;
		Dminus[549] = 12'b000000_000000;
		Dminus[550] = 12'b000000_000000;
		Dminus[551] = 12'b000000_000000;
		Dminus[552] = 12'b000000_000000;
		Dminus[553] = 12'b000000_000000;
		Dminus[554] = 12'b000000_000000;
		Dminus[555] = 12'b000000_000000;
		Dminus[556] = 12'b000000_000000;
		Dminus[557] = 12'b000000_000000;
		Dminus[558] = 12'b000000_000000;
		Dminus[559] = 12'b000000_000000;
		Dminus[560] = 12'b000000_000000;
		Dminus[561] = 12'b000000_000000;
		Dminus[562] = 12'b000000_000000;
		Dminus[563] = 12'b000000_000000;
		Dminus[564] = 12'b000000_000000;
		Dminus[565] = 12'b000000_000000;
		Dminus[566] = 12'b000000_000000;
		Dminus[567] = 12'b000000_000000;
		Dminus[568] = 12'b000000_000000;
		Dminus[569] = 12'b000000_000000;
		Dminus[570] = 12'b000000_000000;
		Dminus[571] = 12'b000000_000000;
		Dminus[572] = 12'b000000_000000;
		Dminus[573] = 12'b000000_000000;
		Dminus[574] = 12'b000000_000000;
		Dminus[575] = 12'b000000_000000;
		Dminus[576] = 12'b000000_000000;
		Dminus[577] = 12'b000000_000000;
		Dminus[578] = 12'b000000_000000;
		Dminus[579] = 12'b000000_000000;
		Dminus[580] = 12'b000000_000000;
		Dminus[581] = 12'b000000_000000;
		Dminus[582] = 12'b000000_000000;
		Dminus[583] = 12'b000000_000000;
		Dminus[584] = 12'b000000_000000;
		Dminus[585] = 12'b000000_000000;
		Dminus[586] = 12'b000000_000000;
		Dminus[587] = 12'b000000_000000;
		Dminus[588] = 12'b000000_000000;
		Dminus[589] = 12'b000000_000000;
		Dminus[590] = 12'b000000_000000;
		Dminus[591] = 12'b000000_000000;
		Dminus[592] = 12'b000000_000000;
		Dminus[593] = 12'b000000_000000;
		Dminus[594] = 12'b000000_000000;
		Dminus[595] = 12'b000000_000000;
		Dminus[596] = 12'b000000_000000;
		Dminus[597] = 12'b000000_000000;
		Dminus[598] = 12'b000000_000000;
		Dminus[599] = 12'b000000_000000;
		Dminus[600] = 12'b000000_000000;
		Dminus[601] = 12'b000000_000000;
		Dminus[602] = 12'b000000_000000;
		Dminus[603] = 12'b000000_000000;
		Dminus[604] = 12'b000000_000000;
		Dminus[605] = 12'b000000_000000;
		Dminus[606] = 12'b000000_000000;
		Dminus[607] = 12'b000000_000000;
		Dminus[608] = 12'b000000_000000;
		Dminus[609] = 12'b000000_000000;
		Dminus[610] = 12'b000000_000000;
		Dminus[611] = 12'b000000_000000;
		Dminus[612] = 12'b000000_000000;
		Dminus[613] = 12'b000000_000000;
		Dminus[614] = 12'b000000_000000;
		Dminus[615] = 12'b000000_000000;
		Dminus[616] = 12'b000000_000000;
		Dminus[617] = 12'b000000_000000;
		Dminus[618] = 12'b000000_000000;
		Dminus[619] = 12'b000000_000000;
		Dminus[620] = 12'b000000_000000;
		Dminus[621] = 12'b000000_000000;
		Dminus[622] = 12'b000000_000000;
		Dminus[623] = 12'b000000_000000;
		Dminus[624] = 12'b000000_000000;
		Dminus[625] = 12'b000000_000000;
		Dminus[626] = 12'b000000_000000;
		Dminus[627] = 12'b000000_000000;
		Dminus[628] = 12'b000000_000000;
		Dminus[629] = 12'b000000_000000;
		Dminus[630] = 12'b000000_000000;
		Dminus[631] = 12'b000000_000000;
		Dminus[632] = 12'b000000_000000;
		Dminus[633] = 12'b000000_000000;
		Dminus[634] = 12'b000000_000000;
		Dminus[635] = 12'b000000_000000;
		Dminus[636] = 12'b000000_000000;
		Dminus[637] = 12'b000000_000000;
		Dminus[638] = 12'b000000_000000;
		Dminus[639] = 12'b000000_000000;
		Dminus[640] = 12'b000000_000000;
		Dminus[641] = 12'b000000_000000;
		Dminus[642] = 12'b000000_000000;
		Dminus[643] = 12'b000000_000000;
		Dminus[644] = 12'b000000_000000;
		Dminus[645] = 12'b000000_000000;
		Dminus[646] = 12'b000000_000000;
		Dminus[647] = 12'b000000_000000;
		Dminus[648] = 12'b000000_000000;
		Dminus[649] = 12'b000000_000000;
		Dminus[650] = 12'b000000_000000;
		Dminus[651] = 12'b000000_000000;
		Dminus[652] = 12'b000000_000000;
		Dminus[653] = 12'b000000_000000;
		Dminus[654] = 12'b000000_000000;
		Dminus[655] = 12'b000000_000000;
		Dminus[656] = 12'b000000_000000;
		Dminus[657] = 12'b000000_000000;
		Dminus[658] = 12'b000000_000000;
		Dminus[659] = 12'b000000_000000;
		Dminus[660] = 12'b000000_000000;
		Dminus[661] = 12'b000000_000000;
		Dminus[662] = 12'b000000_000000;
		Dminus[663] = 12'b000000_000000;
		Dminus[664] = 12'b000000_000000;
		Dminus[665] = 12'b000000_000000;
		Dminus[666] = 12'b000000_000000;
		Dminus[667] = 12'b000000_000000;
		Dminus[668] = 12'b000000_000000;
		Dminus[669] = 12'b000000_000000;
		Dminus[670] = 12'b000000_000000;
		Dminus[671] = 12'b000000_000000;
		Dminus[672] = 12'b000000_000000;
		Dminus[673] = 12'b000000_000000;
		Dminus[674] = 12'b000000_000000;
		Dminus[675] = 12'b000000_000000;
		Dminus[676] = 12'b000000_000000;
		Dminus[677] = 12'b000000_000000;
		Dminus[678] = 12'b000000_000000;
		Dminus[679] = 12'b000000_000000;
		Dminus[680] = 12'b000000_000000;
		Dminus[681] = 12'b000000_000000;
		Dminus[682] = 12'b000000_000000;
		Dminus[683] = 12'b000000_000000;
		Dminus[684] = 12'b000000_000000;
		Dminus[685] = 12'b000000_000000;
		Dminus[686] = 12'b000000_000000;
		Dminus[687] = 12'b000000_000000;
		Dminus[688] = 12'b000000_000000;
		Dminus[689] = 12'b000000_000000;
		Dminus[690] = 12'b000000_000000;
		Dminus[691] = 12'b000000_000000;
		Dminus[692] = 12'b000000_000000;
		Dminus[693] = 12'b000000_000000;
		Dminus[694] = 12'b000000_000000;
		Dminus[695] = 12'b000000_000000;
		Dminus[696] = 12'b000000_000000;
		Dminus[697] = 12'b000000_000000;
		Dminus[698] = 12'b000000_000000;
		Dminus[699] = 12'b000000_000000;
		Dminus[700] = 12'b000000_000000;
		Dminus[701] = 12'b000000_000000;
		Dminus[702] = 12'b000000_000000;
		Dminus[703] = 12'b000000_000000;
		Dminus[704] = 12'b000000_000000;
		Dminus[705] = 12'b000000_000000;
		Dminus[706] = 12'b000000_000000;
		Dminus[707] = 12'b000000_000000;
		Dminus[708] = 12'b000000_000000;
		Dminus[709] = 12'b000000_000000;
		Dminus[710] = 12'b000000_000000;
		Dminus[711] = 12'b000000_000000;
		Dminus[712] = 12'b000000_000000;
		Dminus[713] = 12'b000000_000000;
		Dminus[714] = 12'b000000_000000;
		Dminus[715] = 12'b000000_000000;
		Dminus[716] = 12'b000000_000000;
		Dminus[717] = 12'b000000_000000;
		Dminus[718] = 12'b000000_000000;
		Dminus[719] = 12'b000000_000000;
		Dminus[720] = 12'b000000_000000;
		Dminus[721] = 12'b000000_000000;
		Dminus[722] = 12'b000000_000000;
		Dminus[723] = 12'b000000_000000;
		Dminus[724] = 12'b000000_000000;
		Dminus[725] = 12'b000000_000000;
		Dminus[726] = 12'b000000_000000;
		Dminus[727] = 12'b000000_000000;
		Dminus[728] = 12'b000000_000000;
		Dminus[729] = 12'b000000_000000;
		Dminus[730] = 12'b000000_000000;
		Dminus[731] = 12'b000000_000000;
		Dminus[732] = 12'b000000_000000;
		Dminus[733] = 12'b000000_000000;
		Dminus[734] = 12'b000000_000000;
		Dminus[735] = 12'b000000_000000;
		Dminus[736] = 12'b000000_000000;
		Dminus[737] = 12'b000000_000000;
		Dminus[738] = 12'b000000_000000;
		Dminus[739] = 12'b000000_000000;
		Dminus[740] = 12'b000000_000000;
		Dminus[741] = 12'b000000_000000;
		Dminus[742] = 12'b000000_000000;
		Dminus[743] = 12'b000000_000000;
		Dminus[744] = 12'b000000_000000;
		Dminus[745] = 12'b000000_000000;
		Dminus[746] = 12'b000000_000000;
		Dminus[747] = 12'b000000_000000;
		Dminus[748] = 12'b000000_000000;
		Dminus[749] = 12'b000000_000000;
		Dminus[750] = 12'b000000_000000;
		Dminus[751] = 12'b000000_000000;
		Dminus[752] = 12'b000000_000000;
		Dminus[753] = 12'b000000_000000;
		Dminus[754] = 12'b000000_000000;
		Dminus[755] = 12'b000000_000000;
		Dminus[756] = 12'b000000_000000;
		Dminus[757] = 12'b000000_000000;
		Dminus[758] = 12'b000000_000000;
		Dminus[759] = 12'b000000_000000;
		Dminus[760] = 12'b000000_000000;
		Dminus[761] = 12'b000000_000000;
		Dminus[762] = 12'b000000_000000;
		Dminus[763] = 12'b000000_000000;
		Dminus[764] = 12'b000000_000000;
		Dminus[765] = 12'b000000_000000;
		Dminus[766] = 12'b000000_000000;
		Dminus[767] = 12'b000000_000000;
		Dminus[768] = 12'b000000_000000;
		Dminus[769] = 12'b000000_000000;
		Dminus[770] = 12'b000000_000000;
		Dminus[771] = 12'b000000_000000;
		Dminus[772] = 12'b000000_000000;
		Dminus[773] = 12'b000000_000000;
		Dminus[774] = 12'b000000_000000;
		Dminus[775] = 12'b000000_000000;
		Dminus[776] = 12'b000000_000000;
		Dminus[777] = 12'b000000_000000;
		Dminus[778] = 12'b000000_000000;
		Dminus[779] = 12'b000000_000000;
		Dminus[780] = 12'b000000_000000;
		Dminus[781] = 12'b000000_000000;
		Dminus[782] = 12'b000000_000000;
		Dminus[783] = 12'b000000_000000;
		Dminus[784] = 12'b000000_000000;
		Dminus[785] = 12'b000000_000000;
		Dminus[786] = 12'b000000_000000;
		Dminus[787] = 12'b000000_000000;
		Dminus[788] = 12'b000000_000000;
		Dminus[789] = 12'b000000_000000;
		Dminus[790] = 12'b000000_000000;
		Dminus[791] = 12'b000000_000000;
		Dminus[792] = 12'b000000_000000;
		Dminus[793] = 12'b000000_000000;
		Dminus[794] = 12'b000000_000000;
		Dminus[795] = 12'b000000_000000;
		Dminus[796] = 12'b000000_000000;
		Dminus[797] = 12'b000000_000000;
		Dminus[798] = 12'b000000_000000;
		Dminus[799] = 12'b000000_000000;
		Dminus[800] = 12'b000000_000000;
		Dminus[801] = 12'b000000_000000;
		Dminus[802] = 12'b000000_000000;
		Dminus[803] = 12'b000000_000000;
		Dminus[804] = 12'b000000_000000;
		Dminus[805] = 12'b000000_000000;
		Dminus[806] = 12'b000000_000000;
		Dminus[807] = 12'b000000_000000;
		Dminus[808] = 12'b000000_000000;
		Dminus[809] = 12'b000000_000000;
		Dminus[810] = 12'b000000_000000;
		Dminus[811] = 12'b000000_000000;
		Dminus[812] = 12'b000000_000000;
		Dminus[813] = 12'b000000_000000;
		Dminus[814] = 12'b000000_000000;
		Dminus[815] = 12'b000000_000000;
		Dminus[816] = 12'b000000_000000;
		Dminus[817] = 12'b000000_000000;
		Dminus[818] = 12'b000000_000000;
		Dminus[819] = 12'b000000_000000;
		Dminus[820] = 12'b000000_000000;
		Dminus[821] = 12'b000000_000000;
		Dminus[822] = 12'b000000_000000;
		Dminus[823] = 12'b000000_000000;
		Dminus[824] = 12'b000000_000000;
		Dminus[825] = 12'b000000_000000;
		Dminus[826] = 12'b000000_000000;
		Dminus[827] = 12'b000000_000000;
		Dminus[828] = 12'b000000_000000;
		Dminus[829] = 12'b000000_000000;
		Dminus[830] = 12'b000000_000000;
		Dminus[831] = 12'b000000_000000;
		Dminus[832] = 12'b000000_000000;
		Dminus[833] = 12'b000000_000000;
		Dminus[834] = 12'b000000_000000;
		Dminus[835] = 12'b000000_000000;
		Dminus[836] = 12'b000000_000000;
		Dminus[837] = 12'b000000_000000;
		Dminus[838] = 12'b000000_000000;
		Dminus[839] = 12'b000000_000000;
		Dminus[840] = 12'b000000_000000;
		Dminus[841] = 12'b000000_000000;
		Dminus[842] = 12'b000000_000000;
		Dminus[843] = 12'b000000_000000;
		Dminus[844] = 12'b000000_000000;
		Dminus[845] = 12'b000000_000000;
		Dminus[846] = 12'b000000_000000;
		Dminus[847] = 12'b000000_000000;
		Dminus[848] = 12'b000000_000000;
		Dminus[849] = 12'b000000_000000;
		Dminus[850] = 12'b000000_000000;
		Dminus[851] = 12'b000000_000000;
		Dminus[852] = 12'b000000_000000;
		Dminus[853] = 12'b000000_000000;
		Dminus[854] = 12'b000000_000000;
		Dminus[855] = 12'b000000_000000;
		Dminus[856] = 12'b000000_000000;
		Dminus[857] = 12'b000000_000000;
		Dminus[858] = 12'b000000_000000;
		Dminus[859] = 12'b000000_000000;
		Dminus[860] = 12'b000000_000000;
		Dminus[861] = 12'b000000_000000;
		Dminus[862] = 12'b000000_000000;
		Dminus[863] = 12'b000000_000000;
		Dminus[864] = 12'b000000_000000;
		Dminus[865] = 12'b000000_000000;
		Dminus[866] = 12'b000000_000000;
		Dminus[867] = 12'b000000_000000;
		Dminus[868] = 12'b000000_000000;
		Dminus[869] = 12'b000000_000000;
		Dminus[870] = 12'b000000_000000;
		Dminus[871] = 12'b000000_000000;
		Dminus[872] = 12'b000000_000000;
		Dminus[873] = 12'b000000_000000;
		Dminus[874] = 12'b000000_000000;
		Dminus[875] = 12'b000000_000000;
		Dminus[876] = 12'b000000_000000;
		Dminus[877] = 12'b000000_000000;
		Dminus[878] = 12'b000000_000000;
		Dminus[879] = 12'b000000_000000;
		Dminus[880] = 12'b000000_000000;
		Dminus[881] = 12'b000000_000000;
		Dminus[882] = 12'b000000_000000;
		Dminus[883] = 12'b000000_000000;
		Dminus[884] = 12'b000000_000000;
		Dminus[885] = 12'b000000_000000;
		Dminus[886] = 12'b000000_000000;
		Dminus[887] = 12'b000000_000000;
		Dminus[888] = 12'b000000_000000;
		Dminus[889] = 12'b000000_000000;
		Dminus[890] = 12'b000000_000000;
		Dminus[891] = 12'b000000_000000;
		Dminus[892] = 12'b000000_000000;
		Dminus[893] = 12'b000000_000000;
		Dminus[894] = 12'b000000_000000;
		Dminus[895] = 12'b000000_000000;
		Dminus[896] = 12'b000000_000000;
		Dminus[897] = 12'b000000_000000;
		Dminus[898] = 12'b000000_000000;
		Dminus[899] = 12'b000000_000000;
		Dminus[900] = 12'b000000_000000;
		Dminus[901] = 12'b000000_000000;
		Dminus[902] = 12'b000000_000000;
		Dminus[903] = 12'b000000_000000;
		Dminus[904] = 12'b000000_000000;
		Dminus[905] = 12'b000000_000000;
		Dminus[906] = 12'b000000_000000;
		Dminus[907] = 12'b000000_000000;
		Dminus[908] = 12'b000000_000000;
		Dminus[909] = 12'b000000_000000;
		Dminus[910] = 12'b000000_000000;
		Dminus[911] = 12'b000000_000000;
		Dminus[912] = 12'b000000_000000;
		Dminus[913] = 12'b000000_000000;
		Dminus[914] = 12'b000000_000000;
		Dminus[915] = 12'b000000_000000;
		Dminus[916] = 12'b000000_000000;
		Dminus[917] = 12'b000000_000000;
		Dminus[918] = 12'b000000_000000;
		Dminus[919] = 12'b000000_000000;
		Dminus[920] = 12'b000000_000000;
		Dminus[921] = 12'b000000_000000;
		Dminus[922] = 12'b000000_000000;
		Dminus[923] = 12'b000000_000000;
		Dminus[924] = 12'b000000_000000;
		Dminus[925] = 12'b000000_000000;
		Dminus[926] = 12'b000000_000000;
		Dminus[927] = 12'b000000_000000;
		Dminus[928] = 12'b000000_000000;
		Dminus[929] = 12'b000000_000000;
		Dminus[930] = 12'b000000_000000;
		Dminus[931] = 12'b000000_000000;
		Dminus[932] = 12'b000000_000000;
		Dminus[933] = 12'b000000_000000;
		Dminus[934] = 12'b000000_000000;
		Dminus[935] = 12'b000000_000000;
		Dminus[936] = 12'b000000_000000;
		Dminus[937] = 12'b000000_000000;
		Dminus[938] = 12'b000000_000000;
		Dminus[939] = 12'b000000_000000;
		Dminus[940] = 12'b000000_000000;
		Dminus[941] = 12'b000000_000000;
		Dminus[942] = 12'b000000_000000;
		Dminus[943] = 12'b000000_000000;
		Dminus[944] = 12'b000000_000000;
		Dminus[945] = 12'b000000_000000;
		Dminus[946] = 12'b000000_000000;
		Dminus[947] = 12'b000000_000000;
		Dminus[948] = 12'b000000_000000;
		Dminus[949] = 12'b000000_000000;
		Dminus[950] = 12'b000000_000000;
		Dminus[951] = 12'b000000_000000;
		Dminus[952] = 12'b000000_000000;
		Dminus[953] = 12'b000000_000000;
		Dminus[954] = 12'b000000_000000;
		Dminus[955] = 12'b000000_000000;
		Dminus[956] = 12'b000000_000000;
		Dminus[957] = 12'b000000_000000;
		Dminus[958] = 12'b000000_000000;
		Dminus[959] = 12'b000000_000000;
		Dminus[960] = 12'b000000_000000;
		Dminus[961] = 12'b000000_000000;
		Dminus[962] = 12'b000000_000000;
		Dminus[963] = 12'b000000_000000;
		Dminus[964] = 12'b000000_000000;
		Dminus[965] = 12'b000000_000000;
		Dminus[966] = 12'b000000_000000;
		Dminus[967] = 12'b000000_000000;
		Dminus[968] = 12'b000000_000000;
		Dminus[969] = 12'b000000_000000;
		Dminus[970] = 12'b000000_000000;
		Dminus[971] = 12'b000000_000000;
		Dminus[972] = 12'b000000_000000;
		Dminus[973] = 12'b000000_000000;
		Dminus[974] = 12'b000000_000000;
		Dminus[975] = 12'b000000_000000;
		Dminus[976] = 12'b000000_000000;
		Dminus[977] = 12'b000000_000000;
		Dminus[978] = 12'b000000_000000;
		Dminus[979] = 12'b000000_000000;
		Dminus[980] = 12'b000000_000000;
		Dminus[981] = 12'b000000_000000;
		Dminus[982] = 12'b000000_000000;
		Dminus[983] = 12'b000000_000000;
		Dminus[984] = 12'b000000_000000;
		Dminus[985] = 12'b000000_000000;
		Dminus[986] = 12'b000000_000000;
		Dminus[987] = 12'b000000_000000;
		Dminus[988] = 12'b000000_000000;
		Dminus[989] = 12'b000000_000000;
		Dminus[990] = 12'b000000_000000;
		Dminus[991] = 12'b000000_000000;
		Dminus[992] = 12'b000000_000000;
		Dminus[993] = 12'b000000_000000;
		Dminus[994] = 12'b000000_000000;
		Dminus[995] = 12'b000000_000000;
		Dminus[996] = 12'b000000_000000;
		Dminus[997] = 12'b000000_000000;
		Dminus[998] = 12'b000000_000000;
		Dminus[999] = 12'b000000_000000;
		Dminus[1000] = 12'b000000_000000;
		Dminus[1001] = 12'b000000_000000;
		Dminus[1002] = 12'b000000_000000;
		Dminus[1003] = 12'b000000_000000;
		Dminus[1004] = 12'b000000_000000;
		Dminus[1005] = 12'b000000_000000;
		Dminus[1006] = 12'b000000_000000;
		Dminus[1007] = 12'b000000_000000;
		Dminus[1008] = 12'b000000_000000;
		Dminus[1009] = 12'b000000_000000;
		Dminus[1010] = 12'b000000_000000;
		Dminus[1011] = 12'b000000_000000;
		Dminus[1012] = 12'b000000_000000;
		Dminus[1013] = 12'b000000_000000;
		Dminus[1014] = 12'b000000_000000;
		Dminus[1015] = 12'b000000_000000;
		Dminus[1016] = 12'b000000_000000;
		Dminus[1017] = 12'b000000_000000;
		Dminus[1018] = 12'b000000_000000;
		Dminus[1019] = 12'b000000_000000;
		Dminus[1020] = 12'b000000_000000;
		Dminus[1021] = 12'b000000_000000;
		Dminus[1022] = 12'b000000_000000;
		Dminus[1023] = 12'b000000_000000;
		Dminus[1024] = 12'b000000_000000;
		Dminus[1025] = 12'b000000_000000;
		Dminus[1026] = 12'b000000_000000;
		Dminus[1027] = 12'b000000_000000;
		Dminus[1028] = 12'b000000_000000;
		Dminus[1029] = 12'b000000_000000;
		Dminus[1030] = 12'b000000_000000;
		Dminus[1031] = 12'b000000_000000;
		Dminus[1032] = 12'b000000_000000;
		Dminus[1033] = 12'b000000_000000;
		Dminus[1034] = 12'b000000_000000;
		Dminus[1035] = 12'b000000_000000;
		Dminus[1036] = 12'b000000_000000;
		Dminus[1037] = 12'b000000_000000;
		Dminus[1038] = 12'b000000_000000;
		Dminus[1039] = 12'b000000_000000;
		Dminus[1040] = 12'b000000_000000;
		Dminus[1041] = 12'b000000_000000;
		Dminus[1042] = 12'b000000_000000;
		Dminus[1043] = 12'b000000_000000;
		Dminus[1044] = 12'b000000_000000;
		Dminus[1045] = 12'b000000_000000;
		Dminus[1046] = 12'b000000_000000;
		Dminus[1047] = 12'b000000_000000;
		Dminus[1048] = 12'b000000_000000;
		Dminus[1049] = 12'b000000_000000;
		Dminus[1050] = 12'b000000_000000;
		Dminus[1051] = 12'b000000_000000;
		Dminus[1052] = 12'b000000_000000;
		Dminus[1053] = 12'b000000_000000;
		Dminus[1054] = 12'b000000_000000;
		Dminus[1055] = 12'b000000_000000;
		Dminus[1056] = 12'b000000_000000;
		Dminus[1057] = 12'b000000_000000;
		Dminus[1058] = 12'b000000_000000;
		Dminus[1059] = 12'b000000_000000;
		Dminus[1060] = 12'b000000_000000;
		Dminus[1061] = 12'b000000_000000;
		Dminus[1062] = 12'b000000_000000;
		Dminus[1063] = 12'b000000_000000;
		Dminus[1064] = 12'b000000_000000;
		Dminus[1065] = 12'b000000_000000;
		Dminus[1066] = 12'b000000_000000;
		Dminus[1067] = 12'b000000_000000;
		Dminus[1068] = 12'b000000_000000;
		Dminus[1069] = 12'b000000_000000;
		Dminus[1070] = 12'b000000_000000;
		Dminus[1071] = 12'b000000_000000;
		Dminus[1072] = 12'b000000_000000;
		Dminus[1073] = 12'b000000_000000;
		Dminus[1074] = 12'b000000_000000;
		Dminus[1075] = 12'b000000_000000;
		Dminus[1076] = 12'b000000_000000;
		Dminus[1077] = 12'b000000_000000;
		Dminus[1078] = 12'b000000_000000;
		Dminus[1079] = 12'b000000_000000;
		Dminus[1080] = 12'b000000_000000;
		Dminus[1081] = 12'b000000_000000;
		Dminus[1082] = 12'b000000_000000;
		Dminus[1083] = 12'b000000_000000;
		Dminus[1084] = 12'b000000_000000;
		Dminus[1085] = 12'b000000_000000;
		Dminus[1086] = 12'b000000_000000;
		Dminus[1087] = 12'b000000_000000;
		Dminus[1088] = 12'b000000_000000;
		Dminus[1089] = 12'b000000_000000;
		Dminus[1090] = 12'b000000_000000;
		Dminus[1091] = 12'b000000_000000;
		Dminus[1092] = 12'b000000_000000;
		Dminus[1093] = 12'b000000_000000;
		Dminus[1094] = 12'b000000_000000;
		Dminus[1095] = 12'b000000_000000;
		Dminus[1096] = 12'b000000_000000;
		Dminus[1097] = 12'b000000_000000;
		Dminus[1098] = 12'b000000_000000;
		Dminus[1099] = 12'b000000_000000;
		Dminus[1100] = 12'b000000_000000;
		Dminus[1101] = 12'b000000_000000;
		Dminus[1102] = 12'b000000_000000;
		Dminus[1103] = 12'b000000_000000;
		Dminus[1104] = 12'b000000_000000;
		Dminus[1105] = 12'b000000_000000;
		Dminus[1106] = 12'b000000_000000;
		Dminus[1107] = 12'b000000_000000;
		Dminus[1108] = 12'b000000_000000;
		Dminus[1109] = 12'b000000_000000;
		Dminus[1110] = 12'b000000_000000;
		Dminus[1111] = 12'b000000_000000;
		Dminus[1112] = 12'b000000_000000;
		Dminus[1113] = 12'b000000_000000;
		Dminus[1114] = 12'b000000_000000;
		Dminus[1115] = 12'b000000_000000;
		Dminus[1116] = 12'b000000_000000;
		Dminus[1117] = 12'b000000_000000;
		Dminus[1118] = 12'b000000_000000;
		Dminus[1119] = 12'b000000_000000;
		Dminus[1120] = 12'b000000_000000;
		Dminus[1121] = 12'b000000_000000;
		Dminus[1122] = 12'b000000_000000;
		Dminus[1123] = 12'b000000_000000;
		Dminus[1124] = 12'b000000_000000;
		Dminus[1125] = 12'b000000_000000;
		Dminus[1126] = 12'b000000_000000;
		Dminus[1127] = 12'b000000_000000;
		Dminus[1128] = 12'b000000_000000;
		Dminus[1129] = 12'b000000_000000;
		Dminus[1130] = 12'b000000_000000;
		Dminus[1131] = 12'b000000_000000;
		Dminus[1132] = 12'b000000_000000;
		Dminus[1133] = 12'b000000_000000;
		Dminus[1134] = 12'b000000_000000;
		Dminus[1135] = 12'b000000_000000;
		Dminus[1136] = 12'b000000_000000;
		Dminus[1137] = 12'b000000_000000;
		Dminus[1138] = 12'b000000_000000;
		Dminus[1139] = 12'b000000_000000;
		Dminus[1140] = 12'b000000_000000;
		Dminus[1141] = 12'b000000_000000;
		Dminus[1142] = 12'b000000_000000;
		Dminus[1143] = 12'b000000_000000;
		Dminus[1144] = 12'b000000_000000;
		Dminus[1145] = 12'b000000_000000;
		Dminus[1146] = 12'b000000_000000;
		Dminus[1147] = 12'b000000_000000;
		Dminus[1148] = 12'b000000_000000;
		Dminus[1149] = 12'b000000_000000;
		Dminus[1150] = 12'b000000_000000;
		Dminus[1151] = 12'b000000_000000;
		Dminus[1152] = 12'b000000_000000;
		Dminus[1153] = 12'b000000_000000;
		Dminus[1154] = 12'b000000_000000;
		Dminus[1155] = 12'b000000_000000;
		Dminus[1156] = 12'b000000_000000;
		Dminus[1157] = 12'b000000_000000;
		Dminus[1158] = 12'b000000_000000;
		Dminus[1159] = 12'b000000_000000;
		Dminus[1160] = 12'b000000_000000;
		Dminus[1161] = 12'b000000_000000;
		Dminus[1162] = 12'b000000_000000;
		Dminus[1163] = 12'b000000_000000;
		Dminus[1164] = 12'b000000_000000;
		Dminus[1165] = 12'b000000_000000;
		Dminus[1166] = 12'b000000_000000;
		Dminus[1167] = 12'b000000_000000;
		Dminus[1168] = 12'b000000_000000;
		Dminus[1169] = 12'b000000_000000;
		Dminus[1170] = 12'b000000_000000;
		Dminus[1171] = 12'b000000_000000;
		Dminus[1172] = 12'b000000_000000;
		Dminus[1173] = 12'b000000_000000;
		Dminus[1174] = 12'b000000_000000;
		Dminus[1175] = 12'b000000_000000;
		Dminus[1176] = 12'b000000_000000;
		Dminus[1177] = 12'b000000_000000;
		Dminus[1178] = 12'b000000_000000;
		Dminus[1179] = 12'b000000_000000;
		Dminus[1180] = 12'b000000_000000;
		Dminus[1181] = 12'b000000_000000;
		Dminus[1182] = 12'b000000_000000;
		Dminus[1183] = 12'b000000_000000;
		Dminus[1184] = 12'b000000_000000;
		Dminus[1185] = 12'b000000_000000;
		Dminus[1186] = 12'b000000_000000;
		Dminus[1187] = 12'b000000_000000;
		Dminus[1188] = 12'b000000_000000;
		Dminus[1189] = 12'b000000_000000;
		Dminus[1190] = 12'b000000_000000;
		Dminus[1191] = 12'b000000_000000;
		Dminus[1192] = 12'b000000_000000;
		Dminus[1193] = 12'b000000_000000;
		Dminus[1194] = 12'b000000_000000;
		Dminus[1195] = 12'b000000_000000;
		Dminus[1196] = 12'b000000_000000;
		Dminus[1197] = 12'b000000_000000;
		Dminus[1198] = 12'b000000_000000;
		Dminus[1199] = 12'b000000_000000;
		Dminus[1200] = 12'b000000_000000;
		Dminus[1201] = 12'b000000_000000;
		Dminus[1202] = 12'b000000_000000;
		Dminus[1203] = 12'b000000_000000;
		Dminus[1204] = 12'b000000_000000;
		Dminus[1205] = 12'b000000_000000;
		Dminus[1206] = 12'b000000_000000;
		Dminus[1207] = 12'b000000_000000;
		Dminus[1208] = 12'b000000_000000;
		Dminus[1209] = 12'b000000_000000;
		Dminus[1210] = 12'b000000_000000;
		Dminus[1211] = 12'b000000_000000;
		Dminus[1212] = 12'b000000_000000;
		Dminus[1213] = 12'b000000_000000;
		Dminus[1214] = 12'b000000_000000;
		Dminus[1215] = 12'b000000_000000;
		Dminus[1216] = 12'b000000_000000;
		Dminus[1217] = 12'b000000_000000;
		Dminus[1218] = 12'b000000_000000;
		Dminus[1219] = 12'b000000_000000;
		Dminus[1220] = 12'b000000_000000;
		Dminus[1221] = 12'b000000_000000;
		Dminus[1222] = 12'b000000_000000;
		Dminus[1223] = 12'b000000_000000;
		Dminus[1224] = 12'b000000_000000;
		Dminus[1225] = 12'b000000_000000;
		Dminus[1226] = 12'b000000_000000;
		Dminus[1227] = 12'b000000_000000;
		Dminus[1228] = 12'b000000_000000;
		Dminus[1229] = 12'b000000_000000;
		Dminus[1230] = 12'b000000_000000;
		Dminus[1231] = 12'b000000_000000;
		Dminus[1232] = 12'b000000_000000;
		Dminus[1233] = 12'b000000_000000;
		Dminus[1234] = 12'b000000_000000;
		Dminus[1235] = 12'b000000_000000;
		Dminus[1236] = 12'b000000_000000;
		Dminus[1237] = 12'b000000_000000;
		Dminus[1238] = 12'b000000_000000;
		Dminus[1239] = 12'b000000_000000;
		Dminus[1240] = 12'b000000_000000;
		Dminus[1241] = 12'b000000_000000;
		Dminus[1242] = 12'b000000_000000;
		Dminus[1243] = 12'b000000_000000;
		Dminus[1244] = 12'b000000_000000;
		Dminus[1245] = 12'b000000_000000;
		Dminus[1246] = 12'b000000_000000;
		Dminus[1247] = 12'b000000_000000;
		Dminus[1248] = 12'b000000_000000;
		Dminus[1249] = 12'b000000_000000;
		Dminus[1250] = 12'b000000_000000;
		Dminus[1251] = 12'b000000_000000;
		Dminus[1252] = 12'b000000_000000;
		Dminus[1253] = 12'b000000_000000;
		Dminus[1254] = 12'b000000_000000;
		Dminus[1255] = 12'b000000_000000;
		Dminus[1256] = 12'b000000_000000;
		Dminus[1257] = 12'b000000_000000;
		Dminus[1258] = 12'b000000_000000;
		Dminus[1259] = 12'b000000_000000;
		Dminus[1260] = 12'b000000_000000;
		Dminus[1261] = 12'b000000_000000;
		Dminus[1262] = 12'b000000_000000;
		Dminus[1263] = 12'b000000_000000;
		Dminus[1264] = 12'b000000_000000;
		Dminus[1265] = 12'b000000_000000;
		Dminus[1266] = 12'b000000_000000;
		Dminus[1267] = 12'b000000_000000;
		Dminus[1268] = 12'b000000_000000;
		Dminus[1269] = 12'b000000_000000;
		Dminus[1270] = 12'b000000_000000;
		Dminus[1271] = 12'b000000_000000;
		Dminus[1272] = 12'b000000_000000;
		Dminus[1273] = 12'b000000_000000;
		Dminus[1274] = 12'b000000_000000;
		Dminus[1275] = 12'b000000_000000;
		Dminus[1276] = 12'b000000_000000;
		Dminus[1277] = 12'b000000_000000;
		Dminus[1278] = 12'b000000_000000;
		Dminus[1279] = 12'b000000_000000;
		Dminus[1280] = 12'b000000_000000;
		Dminus[1281] = 12'b000000_000000;
		Dminus[1282] = 12'b000000_000000;
		Dminus[1283] = 12'b000000_000000;
		Dminus[1284] = 12'b000000_000000;
		Dminus[1285] = 12'b000000_000000;
		Dminus[1286] = 12'b000000_000000;
		Dminus[1287] = 12'b000000_000000;
		Dminus[1288] = 12'b000000_000000;
		Dminus[1289] = 12'b000000_000000;
		Dminus[1290] = 12'b000000_000000;
		Dminus[1291] = 12'b000000_000000;
		Dminus[1292] = 12'b000000_000000;
		Dminus[1293] = 12'b000000_000000;
		Dminus[1294] = 12'b000000_000000;
		Dminus[1295] = 12'b000000_000000;
		Dminus[1296] = 12'b000000_000000;
		Dminus[1297] = 12'b000000_000000;
		Dminus[1298] = 12'b000000_000000;
		Dminus[1299] = 12'b000000_000000;
		Dminus[1300] = 12'b000000_000000;
		Dminus[1301] = 12'b000000_000000;
		Dminus[1302] = 12'b000000_000000;
		Dminus[1303] = 12'b000000_000000;
		Dminus[1304] = 12'b000000_000000;
		Dminus[1305] = 12'b000000_000000;
		Dminus[1306] = 12'b000000_000000;
		Dminus[1307] = 12'b000000_000000;
		Dminus[1308] = 12'b000000_000000;
		Dminus[1309] = 12'b000000_000000;
		Dminus[1310] = 12'b000000_000000;
		Dminus[1311] = 12'b000000_000000;
		Dminus[1312] = 12'b000000_000000;
		Dminus[1313] = 12'b000000_000000;
		Dminus[1314] = 12'b000000_000000;
		Dminus[1315] = 12'b000000_000000;
		Dminus[1316] = 12'b000000_000000;
		Dminus[1317] = 12'b000000_000000;
		Dminus[1318] = 12'b000000_000000;
		Dminus[1319] = 12'b000000_000000;
		Dminus[1320] = 12'b000000_000000;
		Dminus[1321] = 12'b000000_000000;
		Dminus[1322] = 12'b000000_000000;
		Dminus[1323] = 12'b000000_000000;
		Dminus[1324] = 12'b000000_000000;
		Dminus[1325] = 12'b000000_000000;
		Dminus[1326] = 12'b000000_000000;
		Dminus[1327] = 12'b000000_000000;
		Dminus[1328] = 12'b000000_000000;
		Dminus[1329] = 12'b000000_000000;
		Dminus[1330] = 12'b000000_000000;
		Dminus[1331] = 12'b000000_000000;
		Dminus[1332] = 12'b000000_000000;
		Dminus[1333] = 12'b000000_000000;
		Dminus[1334] = 12'b000000_000000;
		Dminus[1335] = 12'b000000_000000;
		Dminus[1336] = 12'b000000_000000;
		Dminus[1337] = 12'b000000_000000;
		Dminus[1338] = 12'b000000_000000;
		Dminus[1339] = 12'b000000_000000;
		Dminus[1340] = 12'b000000_000000;
		Dminus[1341] = 12'b000000_000000;
		Dminus[1342] = 12'b000000_000000;
		Dminus[1343] = 12'b000000_000000;
		Dminus[1344] = 12'b000000_000000;
		Dminus[1345] = 12'b000000_000000;
		Dminus[1346] = 12'b000000_000000;
		Dminus[1347] = 12'b000000_000000;
		Dminus[1348] = 12'b000000_000000;
		Dminus[1349] = 12'b000000_000000;
		Dminus[1350] = 12'b000000_000000;
		Dminus[1351] = 12'b000000_000000;
		Dminus[1352] = 12'b000000_000000;
		Dminus[1353] = 12'b000000_000000;
		Dminus[1354] = 12'b000000_000000;
		Dminus[1355] = 12'b000000_000000;
		Dminus[1356] = 12'b000000_000000;
		Dminus[1357] = 12'b000000_000000;
		Dminus[1358] = 12'b000000_000000;
		Dminus[1359] = 12'b000000_000000;
		Dminus[1360] = 12'b000000_000000;
		Dminus[1361] = 12'b000000_000000;
		Dminus[1362] = 12'b000000_000000;
		Dminus[1363] = 12'b000000_000000;
		Dminus[1364] = 12'b000000_000000;
		Dminus[1365] = 12'b000000_000000;
		Dminus[1366] = 12'b000000_000000;
		Dminus[1367] = 12'b000000_000000;
		Dminus[1368] = 12'b000000_000000;
		Dminus[1369] = 12'b000000_000000;
		Dminus[1370] = 12'b000000_000000;
		Dminus[1371] = 12'b000000_000000;
		Dminus[1372] = 12'b000000_000000;
		Dminus[1373] = 12'b000000_000000;
		Dminus[1374] = 12'b000000_000000;
		Dminus[1375] = 12'b000000_000000;
		Dminus[1376] = 12'b000000_000000;
		Dminus[1377] = 12'b000000_000000;
		Dminus[1378] = 12'b000000_000000;
		Dminus[1379] = 12'b000000_000000;
		Dminus[1380] = 12'b000000_000000;
		Dminus[1381] = 12'b000000_000000;
		Dminus[1382] = 12'b000000_000000;
		Dminus[1383] = 12'b000000_000000;
		Dminus[1384] = 12'b000000_000000;
		Dminus[1385] = 12'b000000_000000;
		Dminus[1386] = 12'b000000_000000;
		Dminus[1387] = 12'b000000_000000;
		Dminus[1388] = 12'b000000_000000;
		Dminus[1389] = 12'b000000_000000;
		Dminus[1390] = 12'b000000_000000;
		Dminus[1391] = 12'b000000_000000;
		Dminus[1392] = 12'b000000_000000;
		Dminus[1393] = 12'b000000_000000;
		Dminus[1394] = 12'b000000_000000;
		Dminus[1395] = 12'b000000_000000;
		Dminus[1396] = 12'b000000_000000;
		Dminus[1397] = 12'b000000_000000;
		Dminus[1398] = 12'b000000_000000;
		Dminus[1399] = 12'b000000_000000;
		Dminus[1400] = 12'b000000_000000;
		Dminus[1401] = 12'b000000_000000;
		Dminus[1402] = 12'b000000_000000;
		Dminus[1403] = 12'b000000_000000;
		Dminus[1404] = 12'b000000_000000;
		Dminus[1405] = 12'b000000_000000;
		Dminus[1406] = 12'b000000_000000;
		Dminus[1407] = 12'b000000_000000;
		Dminus[1408] = 12'b000000_000000;
		Dminus[1409] = 12'b000000_000000;
		Dminus[1410] = 12'b000000_000000;
		Dminus[1411] = 12'b000000_000000;
		Dminus[1412] = 12'b000000_000000;
		Dminus[1413] = 12'b000000_000000;
		Dminus[1414] = 12'b000000_000000;
		Dminus[1415] = 12'b000000_000000;
		Dminus[1416] = 12'b000000_000000;
		Dminus[1417] = 12'b000000_000000;
		Dminus[1418] = 12'b000000_000000;
		Dminus[1419] = 12'b000000_000000;
		Dminus[1420] = 12'b000000_000000;
		Dminus[1421] = 12'b000000_000000;
		Dminus[1422] = 12'b000000_000000;
		Dminus[1423] = 12'b000000_000000;
		Dminus[1424] = 12'b000000_000000;
		Dminus[1425] = 12'b000000_000000;
		Dminus[1426] = 12'b000000_000000;
		Dminus[1427] = 12'b000000_000000;
		Dminus[1428] = 12'b000000_000000;
		Dminus[1429] = 12'b000000_000000;
		Dminus[1430] = 12'b000000_000000;
		Dminus[1431] = 12'b000000_000000;
		Dminus[1432] = 12'b000000_000000;
		Dminus[1433] = 12'b000000_000000;
		Dminus[1434] = 12'b000000_000000;
		Dminus[1435] = 12'b000000_000000;
		Dminus[1436] = 12'b000000_000000;
		Dminus[1437] = 12'b000000_000000;
		Dminus[1438] = 12'b000000_000000;
		Dminus[1439] = 12'b000000_000000;
		Dminus[1440] = 12'b000000_000000;
		Dminus[1441] = 12'b000000_000000;
		Dminus[1442] = 12'b000000_000000;
		Dminus[1443] = 12'b000000_000000;
		Dminus[1444] = 12'b000000_000000;
		Dminus[1445] = 12'b000000_000000;
		Dminus[1446] = 12'b000000_000000;
		Dminus[1447] = 12'b000000_000000;
		Dminus[1448] = 12'b000000_000000;
		Dminus[1449] = 12'b000000_000000;
		Dminus[1450] = 12'b000000_000000;
		Dminus[1451] = 12'b000000_000000;
		Dminus[1452] = 12'b000000_000000;
		Dminus[1453] = 12'b000000_000000;
		Dminus[1454] = 12'b000000_000000;
		Dminus[1455] = 12'b000000_000000;
		Dminus[1456] = 12'b000000_000000;
		Dminus[1457] = 12'b000000_000000;
		Dminus[1458] = 12'b000000_000000;
		Dminus[1459] = 12'b000000_000000;
		Dminus[1460] = 12'b000000_000000;
		Dminus[1461] = 12'b000000_000000;
		Dminus[1462] = 12'b000000_000000;
		Dminus[1463] = 12'b000000_000000;
		Dminus[1464] = 12'b000000_000000;
		Dminus[1465] = 12'b000000_000000;
		Dminus[1466] = 12'b000000_000000;
		Dminus[1467] = 12'b000000_000000;
		Dminus[1468] = 12'b000000_000000;
		Dminus[1469] = 12'b000000_000000;
		Dminus[1470] = 12'b000000_000000;
		Dminus[1471] = 12'b000000_000000;
		Dminus[1472] = 12'b000000_000000;
		Dminus[1473] = 12'b000000_000000;
		Dminus[1474] = 12'b000000_000000;
		Dminus[1475] = 12'b000000_000000;
		Dminus[1476] = 12'b000000_000000;
		Dminus[1477] = 12'b000000_000000;
		Dminus[1478] = 12'b000000_000000;
		Dminus[1479] = 12'b000000_000000;
		Dminus[1480] = 12'b000000_000000;
		Dminus[1481] = 12'b000000_000000;
		Dminus[1482] = 12'b000000_000000;
		Dminus[1483] = 12'b000000_000000;
		Dminus[1484] = 12'b000000_000000;
		Dminus[1485] = 12'b000000_000000;
		Dminus[1486] = 12'b000000_000000;
		Dminus[1487] = 12'b000000_000000;
		Dminus[1488] = 12'b000000_000000;
		Dminus[1489] = 12'b000000_000000;
		Dminus[1490] = 12'b000000_000000;
		Dminus[1491] = 12'b000000_000000;
		Dminus[1492] = 12'b000000_000000;
		Dminus[1493] = 12'b000000_000000;
		Dminus[1494] = 12'b000000_000000;
		Dminus[1495] = 12'b000000_000000;
		Dminus[1496] = 12'b000000_000000;
		Dminus[1497] = 12'b000000_000000;
		Dminus[1498] = 12'b000000_000000;
		Dminus[1499] = 12'b000000_000000;
		Dminus[1500] = 12'b000000_000000;
		Dminus[1501] = 12'b000000_000000;
		Dminus[1502] = 12'b000000_000000;
		Dminus[1503] = 12'b000000_000000;
		Dminus[1504] = 12'b000000_000000;
		Dminus[1505] = 12'b000000_000000;
		Dminus[1506] = 12'b000000_000000;
		Dminus[1507] = 12'b000000_000000;
		Dminus[1508] = 12'b000000_000000;
		Dminus[1509] = 12'b000000_000000;
		Dminus[1510] = 12'b000000_000000;
		Dminus[1511] = 12'b000000_000000;
		Dminus[1512] = 12'b000000_000000;
		Dminus[1513] = 12'b000000_000000;
		Dminus[1514] = 12'b000000_000000;
		Dminus[1515] = 12'b000000_000000;
		Dminus[1516] = 12'b000000_000000;
		Dminus[1517] = 12'b000000_000000;
		Dminus[1518] = 12'b000000_000000;
		Dminus[1519] = 12'b000000_000000;
		Dminus[1520] = 12'b000000_000000;
		Dminus[1521] = 12'b000000_000000;
		Dminus[1522] = 12'b000000_000000;
		Dminus[1523] = 12'b000000_000000;
		Dminus[1524] = 12'b000000_000000;
		Dminus[1525] = 12'b000000_000000;
		Dminus[1526] = 12'b000000_000000;
		Dminus[1527] = 12'b000000_000000;
		Dminus[1528] = 12'b000000_000000;
		Dminus[1529] = 12'b000000_000000;
		Dminus[1530] = 12'b000000_000000;
		Dminus[1531] = 12'b000000_000000;
		Dminus[1532] = 12'b000000_000000;
		Dminus[1533] = 12'b000000_000000;
		Dminus[1534] = 12'b000000_000000;
		Dminus[1535] = 12'b000000_000000;
		Dminus[1536] = 12'b000000_000000;
		Dminus[1537] = 12'b000000_000000;
		Dminus[1538] = 12'b000000_000000;
		Dminus[1539] = 12'b000000_000000;
		Dminus[1540] = 12'b000000_000000;
		Dminus[1541] = 12'b000000_000000;
		Dminus[1542] = 12'b000000_000000;
		Dminus[1543] = 12'b000000_000000;
		Dminus[1544] = 12'b000000_000000;
		Dminus[1545] = 12'b000000_000000;
		Dminus[1546] = 12'b000000_000000;
		Dminus[1547] = 12'b000000_000000;
		Dminus[1548] = 12'b000000_000000;
		Dminus[1549] = 12'b000000_000000;
		Dminus[1550] = 12'b000000_000000;
		Dminus[1551] = 12'b000000_000000;
		Dminus[1552] = 12'b000000_000000;
		Dminus[1553] = 12'b000000_000000;
		Dminus[1554] = 12'b000000_000000;
		Dminus[1555] = 12'b000000_000000;
		Dminus[1556] = 12'b000000_000000;
		Dminus[1557] = 12'b000000_000000;
		Dminus[1558] = 12'b000000_000000;
		Dminus[1559] = 12'b000000_000000;
		Dminus[1560] = 12'b000000_000000;
		Dminus[1561] = 12'b000000_000000;
		Dminus[1562] = 12'b000000_000000;
		Dminus[1563] = 12'b000000_000000;
		Dminus[1564] = 12'b000000_000000;
		Dminus[1565] = 12'b000000_000000;
		Dminus[1566] = 12'b000000_000000;
		Dminus[1567] = 12'b000000_000000;
		Dminus[1568] = 12'b000000_000000;
		Dminus[1569] = 12'b000000_000000;
		Dminus[1570] = 12'b000000_000000;
		Dminus[1571] = 12'b000000_000000;
		Dminus[1572] = 12'b000000_000000;
		Dminus[1573] = 12'b000000_000000;
		Dminus[1574] = 12'b000000_000000;
		Dminus[1575] = 12'b000000_000000;
		Dminus[1576] = 12'b000000_000000;
		Dminus[1577] = 12'b000000_000000;
		Dminus[1578] = 12'b000000_000000;
		Dminus[1579] = 12'b000000_000000;
		Dminus[1580] = 12'b000000_000000;
		Dminus[1581] = 12'b000000_000000;
		Dminus[1582] = 12'b000000_000000;
		Dminus[1583] = 12'b000000_000000;
		Dminus[1584] = 12'b000000_000000;
		Dminus[1585] = 12'b000000_000000;
		Dminus[1586] = 12'b000000_000000;
		Dminus[1587] = 12'b000000_000000;
		Dminus[1588] = 12'b000000_000000;
		Dminus[1589] = 12'b000000_000000;
		Dminus[1590] = 12'b000000_000000;
		Dminus[1591] = 12'b000000_000000;
		Dminus[1592] = 12'b000000_000000;
		Dminus[1593] = 12'b000000_000000;
		Dminus[1594] = 12'b000000_000000;
		Dminus[1595] = 12'b000000_000000;
		Dminus[1596] = 12'b000000_000000;
		Dminus[1597] = 12'b000000_000000;
		Dminus[1598] = 12'b000000_000000;
		Dminus[1599] = 12'b000000_000000;
		Dminus[1600] = 12'b000000_000000;
		Dminus[1601] = 12'b000000_000000;
		Dminus[1602] = 12'b000000_000000;
		Dminus[1603] = 12'b000000_000000;
		Dminus[1604] = 12'b000000_000000;
		Dminus[1605] = 12'b000000_000000;
		Dminus[1606] = 12'b000000_000000;
		Dminus[1607] = 12'b000000_000000;
		Dminus[1608] = 12'b000000_000000;
		Dminus[1609] = 12'b000000_000000;
		Dminus[1610] = 12'b000000_000000;
		Dminus[1611] = 12'b000000_000000;
		Dminus[1612] = 12'b000000_000000;
		Dminus[1613] = 12'b000000_000000;
		Dminus[1614] = 12'b000000_000000;
		Dminus[1615] = 12'b000000_000000;
		Dminus[1616] = 12'b000000_000000;
		Dminus[1617] = 12'b000000_000000;
		Dminus[1618] = 12'b000000_000000;
		Dminus[1619] = 12'b000000_000000;
		Dminus[1620] = 12'b000000_000000;
		Dminus[1621] = 12'b000000_000000;
		Dminus[1622] = 12'b000000_000000;
		Dminus[1623] = 12'b000000_000000;
		Dminus[1624] = 12'b000000_000000;
		Dminus[1625] = 12'b000000_000000;
		Dminus[1626] = 12'b000000_000000;
		Dminus[1627] = 12'b000000_000000;
		Dminus[1628] = 12'b000000_000000;
		Dminus[1629] = 12'b000000_000000;
		Dminus[1630] = 12'b000000_000000;
		Dminus[1631] = 12'b000000_000000;
		Dminus[1632] = 12'b000000_000000;
		Dminus[1633] = 12'b000000_000000;
		Dminus[1634] = 12'b000000_000000;
		Dminus[1635] = 12'b000000_000000;
		Dminus[1636] = 12'b000000_000000;
		Dminus[1637] = 12'b000000_000000;
		Dminus[1638] = 12'b000000_000000;
		Dminus[1639] = 12'b000000_000000;
		Dminus[1640] = 12'b000000_000000;
		Dminus[1641] = 12'b000000_000000;
		Dminus[1642] = 12'b000000_000000;
		Dminus[1643] = 12'b000000_000000;
		Dminus[1644] = 12'b000000_000000;
		Dminus[1645] = 12'b000000_000000;
		Dminus[1646] = 12'b000000_000000;
		Dminus[1647] = 12'b000000_000000;
		Dminus[1648] = 12'b000000_000000;
		Dminus[1649] = 12'b000000_000000;
		Dminus[1650] = 12'b000000_000000;
		Dminus[1651] = 12'b000000_000000;
		Dminus[1652] = 12'b000000_000000;
		Dminus[1653] = 12'b000000_000000;
		Dminus[1654] = 12'b000000_000000;
		Dminus[1655] = 12'b000000_000000;
		Dminus[1656] = 12'b000000_000000;
		Dminus[1657] = 12'b000000_000000;
		Dminus[1658] = 12'b000000_000000;
		Dminus[1659] = 12'b000000_000000;
		Dminus[1660] = 12'b000000_000000;
		Dminus[1661] = 12'b000000_000000;
		Dminus[1662] = 12'b000000_000000;
		Dminus[1663] = 12'b000000_000000;
		Dminus[1664] = 12'b000000_000000;
		Dminus[1665] = 12'b000000_000000;
		Dminus[1666] = 12'b000000_000000;
		Dminus[1667] = 12'b000000_000000;
		Dminus[1668] = 12'b000000_000000;
		Dminus[1669] = 12'b000000_000000;
		Dminus[1670] = 12'b000000_000000;
		Dminus[1671] = 12'b000000_000000;
		Dminus[1672] = 12'b000000_000000;
		Dminus[1673] = 12'b000000_000000;
		Dminus[1674] = 12'b000000_000000;
		Dminus[1675] = 12'b000000_000000;
		Dminus[1676] = 12'b000000_000000;
		Dminus[1677] = 12'b000000_000000;
		Dminus[1678] = 12'b000000_000000;
		Dminus[1679] = 12'b000000_000000;
		Dminus[1680] = 12'b000000_000000;
		Dminus[1681] = 12'b000000_000000;
		Dminus[1682] = 12'b000000_000000;
		Dminus[1683] = 12'b000000_000000;
		Dminus[1684] = 12'b000000_000000;
		Dminus[1685] = 12'b000000_000000;
		Dminus[1686] = 12'b000000_000000;
		Dminus[1687] = 12'b000000_000000;
		Dminus[1688] = 12'b000000_000000;
		Dminus[1689] = 12'b000000_000000;
		Dminus[1690] = 12'b000000_000000;
		Dminus[1691] = 12'b000000_000000;
		Dminus[1692] = 12'b000000_000000;
		Dminus[1693] = 12'b000000_000000;
		Dminus[1694] = 12'b000000_000000;
		Dminus[1695] = 12'b000000_000000;
		Dminus[1696] = 12'b000000_000000;
		Dminus[1697] = 12'b000000_000000;
		Dminus[1698] = 12'b000000_000000;
		Dminus[1699] = 12'b000000_000000;
		Dminus[1700] = 12'b000000_000000;
		Dminus[1701] = 12'b000000_000000;
		Dminus[1702] = 12'b000000_000000;
		Dminus[1703] = 12'b000000_000000;
		Dminus[1704] = 12'b000000_000000;
		Dminus[1705] = 12'b000000_000000;
		Dminus[1706] = 12'b000000_000000;
		Dminus[1707] = 12'b000000_000000;
		Dminus[1708] = 12'b000000_000000;
		Dminus[1709] = 12'b000000_000000;
		Dminus[1710] = 12'b000000_000000;
		Dminus[1711] = 12'b000000_000000;
		Dminus[1712] = 12'b000000_000000;
		Dminus[1713] = 12'b000000_000000;
		Dminus[1714] = 12'b000000_000000;
		Dminus[1715] = 12'b000000_000000;
		Dminus[1716] = 12'b000000_000000;
		Dminus[1717] = 12'b000000_000000;
		Dminus[1718] = 12'b000000_000000;
		Dminus[1719] = 12'b000000_000000;
		Dminus[1720] = 12'b000000_000000;
		Dminus[1721] = 12'b000000_000000;
		Dminus[1722] = 12'b000000_000000;
		Dminus[1723] = 12'b000000_000000;
		Dminus[1724] = 12'b000000_000000;
		Dminus[1725] = 12'b000000_000000;
		Dminus[1726] = 12'b000000_000000;
		Dminus[1727] = 12'b000000_000000;
		Dminus[1728] = 12'b000000_000000;
		Dminus[1729] = 12'b000000_000000;
		Dminus[1730] = 12'b000000_000000;
		Dminus[1731] = 12'b000000_000000;
		Dminus[1732] = 12'b000000_000000;
		Dminus[1733] = 12'b000000_000000;
		Dminus[1734] = 12'b000000_000000;
		Dminus[1735] = 12'b000000_000000;
		Dminus[1736] = 12'b000000_000000;
		Dminus[1737] = 12'b000000_000000;
		Dminus[1738] = 12'b000000_000000;
		Dminus[1739] = 12'b000000_000000;
		Dminus[1740] = 12'b000000_000000;
		Dminus[1741] = 12'b000000_000000;
		Dminus[1742] = 12'b000000_000000;
		Dminus[1743] = 12'b000000_000000;
		Dminus[1744] = 12'b000000_000000;
		Dminus[1745] = 12'b000000_000000;
		Dminus[1746] = 12'b000000_000000;
		Dminus[1747] = 12'b000000_000000;
		Dminus[1748] = 12'b000000_000000;
		Dminus[1749] = 12'b000000_000000;
		Dminus[1750] = 12'b000000_000000;
		Dminus[1751] = 12'b000000_000000;
		Dminus[1752] = 12'b000000_000000;
		Dminus[1753] = 12'b000000_000000;
		Dminus[1754] = 12'b000000_000000;
		Dminus[1755] = 12'b000000_000000;
		Dminus[1756] = 12'b000000_000000;
		Dminus[1757] = 12'b000000_000000;
		Dminus[1758] = 12'b000000_000000;
		Dminus[1759] = 12'b000000_000000;
		Dminus[1760] = 12'b000000_000000;
		Dminus[1761] = 12'b000000_000000;
		Dminus[1762] = 12'b000000_000000;
		Dminus[1763] = 12'b000000_000000;
		Dminus[1764] = 12'b000000_000000;
		Dminus[1765] = 12'b000000_000000;
		Dminus[1766] = 12'b000000_000000;
		Dminus[1767] = 12'b000000_000000;
		Dminus[1768] = 12'b000000_000000;
		Dminus[1769] = 12'b000000_000000;
		Dminus[1770] = 12'b000000_000000;
		Dminus[1771] = 12'b000000_000000;
		Dminus[1772] = 12'b000000_000000;
		Dminus[1773] = 12'b000000_000000;
		Dminus[1774] = 12'b000000_000000;
		Dminus[1775] = 12'b000000_000000;
		Dminus[1776] = 12'b000000_000000;
		Dminus[1777] = 12'b000000_000000;
		Dminus[1778] = 12'b000000_000000;
		Dminus[1779] = 12'b000000_000000;
		Dminus[1780] = 12'b000000_000000;
		Dminus[1781] = 12'b000000_000000;
		Dminus[1782] = 12'b000000_000000;
		Dminus[1783] = 12'b000000_000000;
		Dminus[1784] = 12'b000000_000000;
		Dminus[1785] = 12'b000000_000000;
		Dminus[1786] = 12'b000000_000000;
		Dminus[1787] = 12'b000000_000000;
		Dminus[1788] = 12'b000000_000000;
		Dminus[1789] = 12'b000000_000000;
		Dminus[1790] = 12'b000000_000000;
		Dminus[1791] = 12'b000000_000000;
		Dminus[1792] = 12'b000000_000000;
		Dminus[1793] = 12'b000000_000000;
		Dminus[1794] = 12'b000000_000000;
		Dminus[1795] = 12'b000000_000000;
		Dminus[1796] = 12'b000000_000000;
		Dminus[1797] = 12'b000000_000000;
		Dminus[1798] = 12'b000000_000000;
		Dminus[1799] = 12'b000000_000000;
		Dminus[1800] = 12'b000000_000000;
		Dminus[1801] = 12'b000000_000000;
		Dminus[1802] = 12'b000000_000000;
		Dminus[1803] = 12'b000000_000000;
		Dminus[1804] = 12'b000000_000000;
		Dminus[1805] = 12'b000000_000000;
		Dminus[1806] = 12'b000000_000000;
		Dminus[1807] = 12'b000000_000000;
		Dminus[1808] = 12'b000000_000000;
		Dminus[1809] = 12'b000000_000000;
		Dminus[1810] = 12'b000000_000000;
		Dminus[1811] = 12'b000000_000000;
		Dminus[1812] = 12'b000000_000000;
		Dminus[1813] = 12'b000000_000000;
		Dminus[1814] = 12'b000000_000000;
		Dminus[1815] = 12'b000000_000000;
		Dminus[1816] = 12'b000000_000000;
		Dminus[1817] = 12'b000000_000000;
		Dminus[1818] = 12'b000000_000000;
		Dminus[1819] = 12'b000000_000000;
		Dminus[1820] = 12'b000000_000000;
		Dminus[1821] = 12'b000000_000000;
		Dminus[1822] = 12'b000000_000000;
		Dminus[1823] = 12'b000000_000000;
		Dminus[1824] = 12'b000000_000000;
		Dminus[1825] = 12'b000000_000000;
		Dminus[1826] = 12'b000000_000000;
		Dminus[1827] = 12'b000000_000000;
		Dminus[1828] = 12'b000000_000000;
		Dminus[1829] = 12'b000000_000000;
		Dminus[1830] = 12'b000000_000000;
		Dminus[1831] = 12'b000000_000000;
		Dminus[1832] = 12'b000000_000000;
		Dminus[1833] = 12'b000000_000000;
		Dminus[1834] = 12'b000000_000000;
		Dminus[1835] = 12'b000000_000000;
		Dminus[1836] = 12'b000000_000000;
		Dminus[1837] = 12'b000000_000000;
		Dminus[1838] = 12'b000000_000000;
		Dminus[1839] = 12'b000000_000000;
		Dminus[1840] = 12'b000000_000000;
		Dminus[1841] = 12'b000000_000000;
		Dminus[1842] = 12'b000000_000000;
		Dminus[1843] = 12'b000000_000000;
		Dminus[1844] = 12'b000000_000000;
		Dminus[1845] = 12'b000000_000000;
		Dminus[1846] = 12'b000000_000000;
		Dminus[1847] = 12'b000000_000000;
		Dminus[1848] = 12'b000000_000000;
		Dminus[1849] = 12'b000000_000000;
		Dminus[1850] = 12'b000000_000000;
		Dminus[1851] = 12'b000000_000000;
		Dminus[1852] = 12'b000000_000000;
		Dminus[1853] = 12'b000000_000000;
		Dminus[1854] = 12'b000000_000000;
		Dminus[1855] = 12'b000000_000000;
		Dminus[1856] = 12'b000000_000000;
		Dminus[1857] = 12'b000000_000000;
		Dminus[1858] = 12'b000000_000000;
		Dminus[1859] = 12'b000000_000000;
		Dminus[1860] = 12'b000000_000000;
		Dminus[1861] = 12'b000000_000000;
		Dminus[1862] = 12'b000000_000000;
		Dminus[1863] = 12'b000000_000000;
		Dminus[1864] = 12'b000000_000000;
		Dminus[1865] = 12'b000000_000000;
		Dminus[1866] = 12'b000000_000000;
		Dminus[1867] = 12'b000000_000000;
		Dminus[1868] = 12'b000000_000000;
		Dminus[1869] = 12'b000000_000000;
		Dminus[1870] = 12'b000000_000000;
		Dminus[1871] = 12'b000000_000000;
		Dminus[1872] = 12'b000000_000000;
		Dminus[1873] = 12'b000000_000000;
		Dminus[1874] = 12'b000000_000000;
		Dminus[1875] = 12'b000000_000000;
		Dminus[1876] = 12'b000000_000000;
		Dminus[1877] = 12'b000000_000000;
		Dminus[1878] = 12'b000000_000000;
		Dminus[1879] = 12'b000000_000000;
		Dminus[1880] = 12'b000000_000000;
		Dminus[1881] = 12'b000000_000000;
		Dminus[1882] = 12'b000000_000000;
		Dminus[1883] = 12'b000000_000000;
		Dminus[1884] = 12'b000000_000000;
		Dminus[1885] = 12'b000000_000000;
		Dminus[1886] = 12'b000000_000000;
		Dminus[1887] = 12'b000000_000000;
		Dminus[1888] = 12'b000000_000000;
		Dminus[1889] = 12'b000000_000000;
		Dminus[1890] = 12'b000000_000000;
		Dminus[1891] = 12'b000000_000000;
		Dminus[1892] = 12'b000000_000000;
		Dminus[1893] = 12'b000000_000000;
		Dminus[1894] = 12'b000000_000000;
		Dminus[1895] = 12'b000000_000000;
		Dminus[1896] = 12'b000000_000000;
		Dminus[1897] = 12'b000000_000000;
		Dminus[1898] = 12'b000000_000000;
		Dminus[1899] = 12'b000000_000000;
		Dminus[1900] = 12'b000000_000000;
		Dminus[1901] = 12'b000000_000000;
		Dminus[1902] = 12'b000000_000000;
		Dminus[1903] = 12'b000000_000000;
		Dminus[1904] = 12'b000000_000000;
		Dminus[1905] = 12'b000000_000000;
		Dminus[1906] = 12'b000000_000000;
		Dminus[1907] = 12'b000000_000000;
		Dminus[1908] = 12'b000000_000000;
		Dminus[1909] = 12'b000000_000000;
		Dminus[1910] = 12'b000000_000000;
		Dminus[1911] = 12'b000000_000000;
		Dminus[1912] = 12'b000000_000000;
		Dminus[1913] = 12'b000000_000000;
		Dminus[1914] = 12'b000000_000000;
		Dminus[1915] = 12'b000000_000000;
		Dminus[1916] = 12'b000000_000000;
		Dminus[1917] = 12'b000000_000000;
		Dminus[1918] = 12'b000000_000000;
		Dminus[1919] = 12'b000000_000000;
		Dminus[1920] = 12'b000000_000000;
		Dminus[1921] = 12'b000000_000000;
		Dminus[1922] = 12'b000000_000000;
		Dminus[1923] = 12'b000000_000000;
		Dminus[1924] = 12'b000000_000000;
		Dminus[1925] = 12'b000000_000000;
		Dminus[1926] = 12'b000000_000000;
		Dminus[1927] = 12'b000000_000000;
		Dminus[1928] = 12'b000000_000000;
		Dminus[1929] = 12'b000000_000000;
		Dminus[1930] = 12'b000000_000000;
		Dminus[1931] = 12'b000000_000000;
		Dminus[1932] = 12'b000000_000000;
		Dminus[1933] = 12'b000000_000000;
		Dminus[1934] = 12'b000000_000000;
		Dminus[1935] = 12'b000000_000000;
		Dminus[1936] = 12'b000000_000000;
		Dminus[1937] = 12'b000000_000000;
		Dminus[1938] = 12'b000000_000000;
		Dminus[1939] = 12'b000000_000000;
		Dminus[1940] = 12'b000000_000000;
		Dminus[1941] = 12'b000000_000000;
		Dminus[1942] = 12'b000000_000000;
		Dminus[1943] = 12'b000000_000000;
		Dminus[1944] = 12'b000000_000000;
		Dminus[1945] = 12'b000000_000000;
		Dminus[1946] = 12'b000000_000000;
		Dminus[1947] = 12'b000000_000000;
		Dminus[1948] = 12'b000000_000000;
		Dminus[1949] = 12'b000000_000000;
		Dminus[1950] = 12'b000000_000000;
		Dminus[1951] = 12'b000000_000000;
		Dminus[1952] = 12'b000000_000000;
		Dminus[1953] = 12'b000000_000000;
		Dminus[1954] = 12'b000000_000000;
		Dminus[1955] = 12'b000000_000000;
		Dminus[1956] = 12'b000000_000000;
		Dminus[1957] = 12'b000000_000000;
		Dminus[1958] = 12'b000000_000000;
		Dminus[1959] = 12'b000000_000000;
		Dminus[1960] = 12'b000000_000000;
		Dminus[1961] = 12'b000000_000000;
		Dminus[1962] = 12'b000000_000000;
		Dminus[1963] = 12'b000000_000000;
		Dminus[1964] = 12'b000000_000000;
		Dminus[1965] = 12'b000000_000000;
		Dminus[1966] = 12'b000000_000000;
		Dminus[1967] = 12'b000000_000000;
		Dminus[1968] = 12'b000000_000000;
		Dminus[1969] = 12'b000000_000000;
		Dminus[1970] = 12'b000000_000000;
		Dminus[1971] = 12'b000000_000000;
		Dminus[1972] = 12'b000000_000000;
		Dminus[1973] = 12'b000000_000000;
		Dminus[1974] = 12'b000000_000000;
		Dminus[1975] = 12'b000000_000000;
		Dminus[1976] = 12'b000000_000000;
		Dminus[1977] = 12'b000000_000000;
		Dminus[1978] = 12'b000000_000000;
		Dminus[1979] = 12'b000000_000000;
		Dminus[1980] = 12'b000000_000000;
		Dminus[1981] = 12'b000000_000000;
		Dminus[1982] = 12'b000000_000000;
		Dminus[1983] = 12'b000000_000000;
		Dminus[1984] = 12'b000000_000000;
		Dminus[1985] = 12'b000000_000000;
		Dminus[1986] = 12'b000000_000000;
		Dminus[1987] = 12'b000000_000000;
		Dminus[1988] = 12'b000000_000000;
		Dminus[1989] = 12'b000000_000000;
		Dminus[1990] = 12'b000000_000000;
		Dminus[1991] = 12'b000000_000000;
		Dminus[1992] = 12'b000000_000000;
		Dminus[1993] = 12'b000000_000000;
		Dminus[1994] = 12'b000000_000000;
		Dminus[1995] = 12'b000000_000000;
		Dminus[1996] = 12'b000000_000000;
		Dminus[1997] = 12'b000000_000000;
		Dminus[1998] = 12'b000000_000000;
		Dminus[1999] = 12'b000000_000000;
		Dminus[2000] = 12'b000000_000000;
		Dminus[2001] = 12'b000000_000000;
		Dminus[2002] = 12'b000000_000000;
		Dminus[2003] = 12'b000000_000000;
		Dminus[2004] = 12'b000000_000000;
		Dminus[2005] = 12'b000000_000000;
		Dminus[2006] = 12'b000000_000000;
		Dminus[2007] = 12'b000000_000000;
		Dminus[2008] = 12'b000000_000000;
		Dminus[2009] = 12'b000000_000000;
		Dminus[2010] = 12'b000000_000000;
		Dminus[2011] = 12'b000000_000000;
		Dminus[2012] = 12'b000000_000000;
		Dminus[2013] = 12'b000000_000000;
		Dminus[2014] = 12'b000000_000000;
		Dminus[2015] = 12'b000000_000000;
		Dminus[2016] = 12'b000000_000000;
		Dminus[2017] = 12'b000000_000000;
		Dminus[2018] = 12'b000000_000000;
		Dminus[2019] = 12'b000000_000000;
		Dminus[2020] = 12'b000000_000000;
		Dminus[2021] = 12'b000000_000000;
		Dminus[2022] = 12'b000000_000000;
		Dminus[2023] = 12'b000000_000000;
		Dminus[2024] = 12'b000000_000000;
		Dminus[2025] = 12'b000000_000000;
		Dminus[2026] = 12'b000000_000000;
		Dminus[2027] = 12'b000000_000000;
		Dminus[2028] = 12'b000000_000000;
		Dminus[2029] = 12'b000000_000000;
		Dminus[2030] = 12'b000000_000000;
		Dminus[2031] = 12'b000000_000000;
		Dminus[2032] = 12'b000000_000000;
		Dminus[2033] = 12'b000000_000000;
		Dminus[2034] = 12'b000000_000000;
		Dminus[2035] = 12'b000000_000000;
		Dminus[2036] = 12'b000000_000000;
		Dminus[2037] = 12'b000000_000000;
		Dminus[2038] = 12'b000000_000000;
		Dminus[2039] = 12'b000000_000000;
		Dminus[2040] = 12'b000000_000000;
		Dminus[2041] = 12'b000000_000000;
		Dminus[2042] = 12'b000000_000000;
		Dminus[2043] = 12'b000000_000000;
		Dminus[2044] = 12'b000000_000000;
		Dminus[2045] = 12'b000000_000000;
		Dminus[2046] = 12'b000000_000000;
		Dminus[2047] = 12'b000000_000000;
		Dplus[1] = 12'b000000_111111;
		Dplus[2] = 12'b000000_111111;
		Dplus[3] = 12'b000000_111110;
		Dplus[4] = 12'b000000_111101;
		Dplus[5] = 12'b000000_111101;
		Dplus[6] = 12'b000000_111100;
		Dplus[7] = 12'b000000_111011;
		Dplus[8] = 12'b000000_111011;
		Dplus[9] = 12'b000000_111010;
		Dplus[10] = 12'b000000_111001;
		Dplus[11] = 12'b000000_111001;
		Dplus[12] = 12'b000000_111000;
		Dplus[13] = 12'b000000_111000;
		Dplus[14] = 12'b000000_110111;
		Dplus[15] = 12'b000000_110110;
		Dplus[16] = 12'b000000_110110;
		Dplus[17] = 12'b000000_110101;
		Dplus[18] = 12'b000000_110101;
		Dplus[19] = 12'b000000_110100;
		Dplus[20] = 12'b000000_110100;
		Dplus[21] = 12'b000000_110011;
		Dplus[22] = 12'b000000_110010;
		Dplus[23] = 12'b000000_110010;
		Dplus[24] = 12'b000000_110001;
		Dplus[25] = 12'b000000_110001;
		Dplus[26] = 12'b000000_110000;
		Dplus[27] = 12'b000000_110000;
		Dplus[28] = 12'b000000_101111;
		Dplus[29] = 12'b000000_101111;
		Dplus[30] = 12'b000000_101110;
		Dplus[31] = 12'b000000_101110;
		Dplus[32] = 12'b000000_101101;
		Dplus[33] = 12'b000000_101101;
		Dplus[34] = 12'b000000_101100;
		Dplus[35] = 12'b000000_101100;
		Dplus[36] = 12'b000000_101011;
		Dplus[37] = 12'b000000_101011;
		Dplus[38] = 12'b000000_101010;
		Dplus[39] = 12'b000000_101010;
		Dplus[40] = 12'b000000_101001;
		Dplus[41] = 12'b000000_101001;
		Dplus[42] = 12'b000000_101001;
		Dplus[43] = 12'b000000_101000;
		Dplus[44] = 12'b000000_101000;
		Dplus[45] = 12'b000000_100111;
		Dplus[46] = 12'b000000_100111;
		Dplus[47] = 12'b000000_100110;
		Dplus[48] = 12'b000000_100110;
		Dplus[49] = 12'b000000_100110;
		Dplus[50] = 12'b000000_100101;
		Dplus[51] = 12'b000000_100101;
		Dplus[52] = 12'b000000_100100;
		Dplus[53] = 12'b000000_100100;
		Dplus[54] = 12'b000000_100100;
		Dplus[55] = 12'b000000_100011;
		Dplus[56] = 12'b000000_100011;
		Dplus[57] = 12'b000000_100011;
		Dplus[58] = 12'b000000_100010;
		Dplus[59] = 12'b000000_100010;
		Dplus[60] = 12'b000000_100001;
		Dplus[61] = 12'b000000_100001;
		Dplus[62] = 12'b000000_100001;
		Dplus[63] = 12'b000000_100000;
		Dplus[64] = 12'b000000_100000;
		Dplus[65] = 12'b000000_100000;
		Dplus[66] = 12'b000000_011111;
		Dplus[67] = 12'b000000_011111;
		Dplus[68] = 12'b000000_011111;
		Dplus[69] = 12'b000000_011110;
		Dplus[70] = 12'b000000_011110;
		Dplus[71] = 12'b000000_011110;
		Dplus[72] = 12'b000000_011101;
		Dplus[73] = 12'b000000_011101;
		Dplus[74] = 12'b000000_011101;
		Dplus[75] = 12'b000000_011100;
		Dplus[76] = 12'b000000_011100;
		Dplus[77] = 12'b000000_011100;
		Dplus[78] = 12'b000000_011011;
		Dplus[79] = 12'b000000_011011;
		Dplus[80] = 12'b000000_011011;
		Dplus[81] = 12'b000000_011011;
		Dplus[82] = 12'b000000_011010;
		Dplus[83] = 12'b000000_011010;
		Dplus[84] = 12'b000000_011010;
		Dplus[85] = 12'b000000_011001;
		Dplus[86] = 12'b000000_011001;
		Dplus[87] = 12'b000000_011001;
		Dplus[88] = 12'b000000_011001;
		Dplus[89] = 12'b000000_011000;
		Dplus[90] = 12'b000000_011000;
		Dplus[91] = 12'b000000_011000;
		Dplus[92] = 12'b000000_011000;
		Dplus[93] = 12'b000000_010111;
		Dplus[94] = 12'b000000_010111;
		Dplus[95] = 12'b000000_010111;
		Dplus[96] = 12'b000000_010111;
		Dplus[97] = 12'b000000_010110;
		Dplus[98] = 12'b000000_010110;
		Dplus[99] = 12'b000000_010110;
		Dplus[100] = 12'b000000_010110;
		Dplus[101] = 12'b000000_010101;
		Dplus[102] = 12'b000000_010101;
		Dplus[103] = 12'b000000_010101;
		Dplus[104] = 12'b000000_010101;
		Dplus[105] = 12'b000000_010101;
		Dplus[106] = 12'b000000_010100;
		Dplus[107] = 12'b000000_010100;
		Dplus[108] = 12'b000000_010100;
		Dplus[109] = 12'b000000_010100;
		Dplus[110] = 12'b000000_010011;
		Dplus[111] = 12'b000000_010011;
		Dplus[112] = 12'b000000_010011;
		Dplus[113] = 12'b000000_010011;
		Dplus[114] = 12'b000000_010011;
		Dplus[115] = 12'b000000_010010;
		Dplus[116] = 12'b000000_010010;
		Dplus[117] = 12'b000000_010010;
		Dplus[118] = 12'b000000_010010;
		Dplus[119] = 12'b000000_010010;
		Dplus[120] = 12'b000000_010001;
		Dplus[121] = 12'b000000_010001;
		Dplus[122] = 12'b000000_010001;
		Dplus[123] = 12'b000000_010001;
		Dplus[124] = 12'b000000_010001;
		Dplus[125] = 12'b000000_010001;
		Dplus[126] = 12'b000000_010000;
		Dplus[127] = 12'b000000_010000;
		Dplus[128] = 12'b000000_010000;
		Dplus[129] = 12'b000000_010000;
		Dplus[130] = 12'b000000_010000;
		Dplus[131] = 12'b000000_001111;
		Dplus[132] = 12'b000000_001111;
		Dplus[133] = 12'b000000_001111;
		Dplus[134] = 12'b000000_001111;
		Dplus[135] = 12'b000000_001111;
		Dplus[136] = 12'b000000_001111;
		Dplus[137] = 12'b000000_001111;
		Dplus[138] = 12'b000000_001110;
		Dplus[139] = 12'b000000_001110;
		Dplus[140] = 12'b000000_001110;
		Dplus[141] = 12'b000000_001110;
		Dplus[142] = 12'b000000_001110;
		Dplus[143] = 12'b000000_001110;
		Dplus[144] = 12'b000000_001101;
		Dplus[145] = 12'b000000_001101;
		Dplus[146] = 12'b000000_001101;
		Dplus[147] = 12'b000000_001101;
		Dplus[148] = 12'b000000_001101;
		Dplus[149] = 12'b000000_001101;
		Dplus[150] = 12'b000000_001101;
		Dplus[151] = 12'b000000_001100;
		Dplus[152] = 12'b000000_001100;
		Dplus[153] = 12'b000000_001100;
		Dplus[154] = 12'b000000_001100;
		Dplus[155] = 12'b000000_001100;
		Dplus[156] = 12'b000000_001100;
		Dplus[157] = 12'b000000_001100;
		Dplus[158] = 12'b000000_001100;
		Dplus[159] = 12'b000000_001011;
		Dplus[160] = 12'b000000_001011;
		Dplus[161] = 12'b000000_001011;
		Dplus[162] = 12'b000000_001011;
		Dplus[163] = 12'b000000_001011;
		Dplus[164] = 12'b000000_001011;
		Dplus[165] = 12'b000000_001011;
		Dplus[166] = 12'b000000_001011;
		Dplus[167] = 12'b000000_001010;
		Dplus[168] = 12'b000000_001010;
		Dplus[169] = 12'b000000_001010;
		Dplus[170] = 12'b000000_001010;
		Dplus[171] = 12'b000000_001010;
		Dplus[172] = 12'b000000_001010;
		Dplus[173] = 12'b000000_001010;
		Dplus[174] = 12'b000000_001010;
		Dplus[175] = 12'b000000_001010;
		Dplus[176] = 12'b000000_001010;
		Dplus[177] = 12'b000000_001001;
		Dplus[178] = 12'b000000_001001;
		Dplus[179] = 12'b000000_001001;
		Dplus[180] = 12'b000000_001001;
		Dplus[181] = 12'b000000_001001;
		Dplus[182] = 12'b000000_001001;
		Dplus[183] = 12'b000000_001001;
		Dplus[184] = 12'b000000_001001;
		Dplus[185] = 12'b000000_001001;
		Dplus[186] = 12'b000000_001001;
		Dplus[187] = 12'b000000_001000;
		Dplus[188] = 12'b000000_001000;
		Dplus[189] = 12'b000000_001000;
		Dplus[190] = 12'b000000_001000;
		Dplus[191] = 12'b000000_001000;
		Dplus[192] = 12'b000000_001000;
		Dplus[193] = 12'b000000_001000;
		Dplus[194] = 12'b000000_001000;
		Dplus[195] = 12'b000000_001000;
		Dplus[196] = 12'b000000_001000;
		Dplus[197] = 12'b000000_001000;
		Dplus[198] = 12'b000000_000111;
		Dplus[199] = 12'b000000_000111;
		Dplus[200] = 12'b000000_000111;
		Dplus[201] = 12'b000000_000111;
		Dplus[202] = 12'b000000_000111;
		Dplus[203] = 12'b000000_000111;
		Dplus[204] = 12'b000000_000111;
		Dplus[205] = 12'b000000_000111;
		Dplus[206] = 12'b000000_000111;
		Dplus[207] = 12'b000000_000111;
		Dplus[208] = 12'b000000_000111;
		Dplus[209] = 12'b000000_000111;
		Dplus[210] = 12'b000000_000111;
		Dplus[211] = 12'b000000_000111;
		Dplus[212] = 12'b000000_000110;
		Dplus[213] = 12'b000000_000110;
		Dplus[214] = 12'b000000_000110;
		Dplus[215] = 12'b000000_000110;
		Dplus[216] = 12'b000000_000110;
		Dplus[217] = 12'b000000_000110;
		Dplus[218] = 12'b000000_000110;
		Dplus[219] = 12'b000000_000110;
		Dplus[220] = 12'b000000_000110;
		Dplus[221] = 12'b000000_000110;
		Dplus[222] = 12'b000000_000110;
		Dplus[223] = 12'b000000_000110;
		Dplus[224] = 12'b000000_000110;
		Dplus[225] = 12'b000000_000110;
		Dplus[226] = 12'b000000_000110;
		Dplus[227] = 12'b000000_000101;
		Dplus[228] = 12'b000000_000101;
		Dplus[229] = 12'b000000_000101;
		Dplus[230] = 12'b000000_000101;
		Dplus[231] = 12'b000000_000101;
		Dplus[232] = 12'b000000_000101;
		Dplus[233] = 12'b000000_000101;
		Dplus[234] = 12'b000000_000101;
		Dplus[235] = 12'b000000_000101;
		Dplus[236] = 12'b000000_000101;
		Dplus[237] = 12'b000000_000101;
		Dplus[238] = 12'b000000_000101;
		Dplus[239] = 12'b000000_000101;
		Dplus[240] = 12'b000000_000101;
		Dplus[241] = 12'b000000_000101;
		Dplus[242] = 12'b000000_000101;
		Dplus[243] = 12'b000000_000101;
		Dplus[244] = 12'b000000_000101;
		Dplus[245] = 12'b000000_000101;
		Dplus[246] = 12'b000000_000100;
		Dplus[247] = 12'b000000_000100;
		Dplus[248] = 12'b000000_000100;
		Dplus[249] = 12'b000000_000100;
		Dplus[250] = 12'b000000_000100;
		Dplus[251] = 12'b000000_000100;
		Dplus[252] = 12'b000000_000100;
		Dplus[253] = 12'b000000_000100;
		Dplus[254] = 12'b000000_000100;
		Dplus[255] = 12'b000000_000100;
		Dplus[256] = 12'b000000_000100;
		Dplus[257] = 12'b000000_000100;
		Dplus[258] = 12'b000000_000100;
		Dplus[259] = 12'b000000_000100;
		Dplus[260] = 12'b000000_000100;
		Dplus[261] = 12'b000000_000100;
		Dplus[262] = 12'b000000_000100;
		Dplus[263] = 12'b000000_000100;
		Dplus[264] = 12'b000000_000100;
		Dplus[265] = 12'b000000_000100;
		Dplus[266] = 12'b000000_000100;
		Dplus[267] = 12'b000000_000100;
		Dplus[268] = 12'b000000_000100;
		Dplus[269] = 12'b000000_000011;
		Dplus[270] = 12'b000000_000011;
		Dplus[271] = 12'b000000_000011;
		Dplus[272] = 12'b000000_000011;
		Dplus[273] = 12'b000000_000011;
		Dplus[274] = 12'b000000_000011;
		Dplus[275] = 12'b000000_000011;
		Dplus[276] = 12'b000000_000011;
		Dplus[277] = 12'b000000_000011;
		Dplus[278] = 12'b000000_000011;
		Dplus[279] = 12'b000000_000011;
		Dplus[280] = 12'b000000_000011;
		Dplus[281] = 12'b000000_000011;
		Dplus[282] = 12'b000000_000011;
		Dplus[283] = 12'b000000_000011;
		Dplus[284] = 12'b000000_000011;
		Dplus[285] = 12'b000000_000011;
		Dplus[286] = 12'b000000_000011;
		Dplus[287] = 12'b000000_000011;
		Dplus[288] = 12'b000000_000011;
		Dplus[289] = 12'b000000_000011;
		Dplus[290] = 12'b000000_000011;
		Dplus[291] = 12'b000000_000011;
		Dplus[292] = 12'b000000_000011;
		Dplus[293] = 12'b000000_000011;
		Dplus[294] = 12'b000000_000011;
		Dplus[295] = 12'b000000_000011;
		Dplus[296] = 12'b000000_000011;
		Dplus[297] = 12'b000000_000011;
		Dplus[298] = 12'b000000_000011;
		Dplus[299] = 12'b000000_000011;
		Dplus[300] = 12'b000000_000010;
		Dplus[301] = 12'b000000_000010;
		Dplus[302] = 12'b000000_000010;
		Dplus[303] = 12'b000000_000010;
		Dplus[304] = 12'b000000_000010;
		Dplus[305] = 12'b000000_000010;
		Dplus[306] = 12'b000000_000010;
		Dplus[307] = 12'b000000_000010;
		Dplus[308] = 12'b000000_000010;
		Dplus[309] = 12'b000000_000010;
		Dplus[310] = 12'b000000_000010;
		Dplus[311] = 12'b000000_000010;
		Dplus[312] = 12'b000000_000010;
		Dplus[313] = 12'b000000_000010;
		Dplus[314] = 12'b000000_000010;
		Dplus[315] = 12'b000000_000010;
		Dplus[316] = 12'b000000_000010;
		Dplus[317] = 12'b000000_000010;
		Dplus[318] = 12'b000000_000010;
		Dplus[319] = 12'b000000_000010;
		Dplus[320] = 12'b000000_000010;
		Dplus[321] = 12'b000000_000010;
		Dplus[322] = 12'b000000_000010;
		Dplus[323] = 12'b000000_000010;
		Dplus[324] = 12'b000000_000010;
		Dplus[325] = 12'b000000_000010;
		Dplus[326] = 12'b000000_000010;
		Dplus[327] = 12'b000000_000010;
		Dplus[328] = 12'b000000_000010;
		Dplus[329] = 12'b000000_000010;
		Dplus[330] = 12'b000000_000010;
		Dplus[331] = 12'b000000_000010;
		Dplus[332] = 12'b000000_000010;
		Dplus[333] = 12'b000000_000010;
		Dplus[334] = 12'b000000_000010;
		Dplus[335] = 12'b000000_000010;
		Dplus[336] = 12'b000000_000010;
		Dplus[337] = 12'b000000_000010;
		Dplus[338] = 12'b000000_000010;
		Dplus[339] = 12'b000000_000010;
		Dplus[340] = 12'b000000_000010;
		Dplus[341] = 12'b000000_000010;
		Dplus[342] = 12'b000000_000010;
		Dplus[343] = 12'b000000_000010;
		Dplus[344] = 12'b000000_000010;
		Dplus[345] = 12'b000000_000010;
		Dplus[346] = 12'b000000_000010;
		Dplus[347] = 12'b000000_000001;
		Dplus[348] = 12'b000000_000001;
		Dplus[349] = 12'b000000_000001;
		Dplus[350] = 12'b000000_000001;
		Dplus[351] = 12'b000000_000001;
		Dplus[352] = 12'b000000_000001;
		Dplus[353] = 12'b000000_000001;
		Dplus[354] = 12'b000000_000001;
		Dplus[355] = 12'b000000_000001;
		Dplus[356] = 12'b000000_000001;
		Dplus[357] = 12'b000000_000001;
		Dplus[358] = 12'b000000_000001;
		Dplus[359] = 12'b000000_000001;
		Dplus[360] = 12'b000000_000001;
		Dplus[361] = 12'b000000_000001;
		Dplus[362] = 12'b000000_000001;
		Dplus[363] = 12'b000000_000001;
		Dplus[364] = 12'b000000_000001;
		Dplus[365] = 12'b000000_000001;
		Dplus[366] = 12'b000000_000001;
		Dplus[367] = 12'b000000_000001;
		Dplus[368] = 12'b000000_000001;
		Dplus[369] = 12'b000000_000001;
		Dplus[370] = 12'b000000_000001;
		Dplus[371] = 12'b000000_000001;
		Dplus[372] = 12'b000000_000001;
		Dplus[373] = 12'b000000_000001;
		Dplus[374] = 12'b000000_000001;
		Dplus[375] = 12'b000000_000001;
		Dplus[376] = 12'b000000_000001;
		Dplus[377] = 12'b000000_000001;
		Dplus[378] = 12'b000000_000001;
		Dplus[379] = 12'b000000_000001;
		Dplus[380] = 12'b000000_000001;
		Dplus[381] = 12'b000000_000001;
		Dplus[382] = 12'b000000_000001;
		Dplus[383] = 12'b000000_000001;
		Dplus[384] = 12'b000000_000001;
		Dplus[385] = 12'b000000_000001;
		Dplus[386] = 12'b000000_000001;
		Dplus[387] = 12'b000000_000001;
		Dplus[388] = 12'b000000_000001;
		Dplus[389] = 12'b000000_000001;
		Dplus[390] = 12'b000000_000001;
		Dplus[391] = 12'b000000_000001;
		Dplus[392] = 12'b000000_000001;
		Dplus[393] = 12'b000000_000001;
		Dplus[394] = 12'b000000_000001;
		Dplus[395] = 12'b000000_000001;
		Dplus[396] = 12'b000000_000001;
		Dplus[397] = 12'b000000_000001;
		Dplus[398] = 12'b000000_000001;
		Dplus[399] = 12'b000000_000001;
		Dplus[400] = 12'b000000_000001;
		Dplus[401] = 12'b000000_000001;
		Dplus[402] = 12'b000000_000001;
		Dplus[403] = 12'b000000_000001;
		Dplus[404] = 12'b000000_000001;
		Dplus[405] = 12'b000000_000001;
		Dplus[406] = 12'b000000_000001;
		Dplus[407] = 12'b000000_000001;
		Dplus[408] = 12'b000000_000001;
		Dplus[409] = 12'b000000_000001;
		Dplus[410] = 12'b000000_000001;
		Dplus[411] = 12'b000000_000001;
		Dplus[412] = 12'b000000_000001;
		Dplus[413] = 12'b000000_000001;
		Dplus[414] = 12'b000000_000001;
		Dplus[415] = 12'b000000_000001;
		Dplus[416] = 12'b000000_000001;
		Dplus[417] = 12'b000000_000001;
		Dplus[418] = 12'b000000_000001;
		Dplus[419] = 12'b000000_000001;
		Dplus[420] = 12'b000000_000001;
		Dplus[421] = 12'b000000_000001;
		Dplus[422] = 12'b000000_000001;
		Dplus[423] = 12'b000000_000001;
		Dplus[424] = 12'b000000_000001;
		Dplus[425] = 12'b000000_000001;
		Dplus[426] = 12'b000000_000001;
		Dplus[427] = 12'b000000_000001;
		Dplus[428] = 12'b000000_000001;
		Dplus[429] = 12'b000000_000001;
		Dplus[430] = 12'b000000_000001;
		Dplus[431] = 12'b000000_000001;
		Dplus[432] = 12'b000000_000001;
		Dplus[433] = 12'b000000_000001;
		Dplus[434] = 12'b000000_000001;
		Dplus[435] = 12'b000000_000001;
		Dplus[436] = 12'b000000_000001;
		Dplus[437] = 12'b000000_000001;
		Dplus[438] = 12'b000000_000001;
		Dplus[439] = 12'b000000_000001;
		Dplus[440] = 12'b000000_000001;
		Dplus[441] = 12'b000000_000001;
		Dplus[442] = 12'b000000_000001;
		Dplus[443] = 12'b000000_000001;
		Dplus[444] = 12'b000000_000001;
		Dplus[445] = 12'b000000_000001;
		Dplus[446] = 12'b000000_000001;
		Dplus[447] = 12'b000000_000001;
		Dplus[448] = 12'b000000_000000;
		Dplus[449] = 12'b000000_000000;
		Dplus[450] = 12'b000000_000000;
		Dplus[451] = 12'b000000_000000;
		Dplus[452] = 12'b000000_000000;
		Dplus[453] = 12'b000000_000000;
		Dplus[454] = 12'b000000_000000;
		Dplus[455] = 12'b000000_000000;
		Dplus[456] = 12'b000000_000000;
		Dplus[457] = 12'b000000_000000;
		Dplus[458] = 12'b000000_000000;
		Dplus[459] = 12'b000000_000000;
		Dplus[460] = 12'b000000_000000;
		Dplus[461] = 12'b000000_000000;
		Dplus[462] = 12'b000000_000000;
		Dplus[463] = 12'b000000_000000;
		Dplus[464] = 12'b000000_000000;
		Dplus[465] = 12'b000000_000000;
		Dplus[466] = 12'b000000_000000;
		Dplus[467] = 12'b000000_000000;
		Dplus[468] = 12'b000000_000000;
		Dplus[469] = 12'b000000_000000;
		Dplus[470] = 12'b000000_000000;
		Dplus[471] = 12'b000000_000000;
		Dplus[472] = 12'b000000_000000;
		Dplus[473] = 12'b000000_000000;
		Dplus[474] = 12'b000000_000000;
		Dplus[475] = 12'b000000_000000;
		Dplus[476] = 12'b000000_000000;
		Dplus[477] = 12'b000000_000000;
		Dplus[478] = 12'b000000_000000;
		Dplus[479] = 12'b000000_000000;
		Dplus[480] = 12'b000000_000000;
		Dplus[481] = 12'b000000_000000;
		Dplus[482] = 12'b000000_000000;
		Dplus[483] = 12'b000000_000000;
		Dplus[484] = 12'b000000_000000;
		Dplus[485] = 12'b000000_000000;
		Dplus[486] = 12'b000000_000000;
		Dplus[487] = 12'b000000_000000;
		Dplus[488] = 12'b000000_000000;
		Dplus[489] = 12'b000000_000000;
		Dplus[490] = 12'b000000_000000;
		Dplus[491] = 12'b000000_000000;
		Dplus[492] = 12'b000000_000000;
		Dplus[493] = 12'b000000_000000;
		Dplus[494] = 12'b000000_000000;
		Dplus[495] = 12'b000000_000000;
		Dplus[496] = 12'b000000_000000;
		Dplus[497] = 12'b000000_000000;
		Dplus[498] = 12'b000000_000000;
		Dplus[499] = 12'b000000_000000;
		Dplus[500] = 12'b000000_000000;
		Dplus[501] = 12'b000000_000000;
		Dplus[502] = 12'b000000_000000;
		Dplus[503] = 12'b000000_000000;
		Dplus[504] = 12'b000000_000000;
		Dplus[505] = 12'b000000_000000;
		Dplus[506] = 12'b000000_000000;
		Dplus[507] = 12'b000000_000000;
		Dplus[508] = 12'b000000_000000;
		Dplus[509] = 12'b000000_000000;
		Dplus[510] = 12'b000000_000000;
		Dplus[511] = 12'b000000_000000;
		Dplus[512] = 12'b000000_000000;
		Dplus[513] = 12'b000000_000000;
		Dplus[514] = 12'b000000_000000;
		Dplus[515] = 12'b000000_000000;
		Dplus[516] = 12'b000000_000000;
		Dplus[517] = 12'b000000_000000;
		Dplus[518] = 12'b000000_000000;
		Dplus[519] = 12'b000000_000000;
		Dplus[520] = 12'b000000_000000;
		Dplus[521] = 12'b000000_000000;
		Dplus[522] = 12'b000000_000000;
		Dplus[523] = 12'b000000_000000;
		Dplus[524] = 12'b000000_000000;
		Dplus[525] = 12'b000000_000000;
		Dplus[526] = 12'b000000_000000;
		Dplus[527] = 12'b000000_000000;
		Dplus[528] = 12'b000000_000000;
		Dplus[529] = 12'b000000_000000;
		Dplus[530] = 12'b000000_000000;
		Dplus[531] = 12'b000000_000000;
		Dplus[532] = 12'b000000_000000;
		Dplus[533] = 12'b000000_000000;
		Dplus[534] = 12'b000000_000000;
		Dplus[535] = 12'b000000_000000;
		Dplus[536] = 12'b000000_000000;
		Dplus[537] = 12'b000000_000000;
		Dplus[538] = 12'b000000_000000;
		Dplus[539] = 12'b000000_000000;
		Dplus[540] = 12'b000000_000000;
		Dplus[541] = 12'b000000_000000;
		Dplus[542] = 12'b000000_000000;
		Dplus[543] = 12'b000000_000000;
		Dplus[544] = 12'b000000_000000;
		Dplus[545] = 12'b000000_000000;
		Dplus[546] = 12'b000000_000000;
		Dplus[547] = 12'b000000_000000;
		Dplus[548] = 12'b000000_000000;
		Dplus[549] = 12'b000000_000000;
		Dplus[550] = 12'b000000_000000;
		Dplus[551] = 12'b000000_000000;
		Dplus[552] = 12'b000000_000000;
		Dplus[553] = 12'b000000_000000;
		Dplus[554] = 12'b000000_000000;
		Dplus[555] = 12'b000000_000000;
		Dplus[556] = 12'b000000_000000;
		Dplus[557] = 12'b000000_000000;
		Dplus[558] = 12'b000000_000000;
		Dplus[559] = 12'b000000_000000;
		Dplus[560] = 12'b000000_000000;
		Dplus[561] = 12'b000000_000000;
		Dplus[562] = 12'b000000_000000;
		Dplus[563] = 12'b000000_000000;
		Dplus[564] = 12'b000000_000000;
		Dplus[565] = 12'b000000_000000;
		Dplus[566] = 12'b000000_000000;
		Dplus[567] = 12'b000000_000000;
		Dplus[568] = 12'b000000_000000;
		Dplus[569] = 12'b000000_000000;
		Dplus[570] = 12'b000000_000000;
		Dplus[571] = 12'b000000_000000;
		Dplus[572] = 12'b000000_000000;
		Dplus[573] = 12'b000000_000000;
		Dplus[574] = 12'b000000_000000;
		Dplus[575] = 12'b000000_000000;
		Dplus[576] = 12'b000000_000000;
		Dplus[577] = 12'b000000_000000;
		Dplus[578] = 12'b000000_000000;
		Dplus[579] = 12'b000000_000000;
		Dplus[580] = 12'b000000_000000;
		Dplus[581] = 12'b000000_000000;
		Dplus[582] = 12'b000000_000000;
		Dplus[583] = 12'b000000_000000;
		Dplus[584] = 12'b000000_000000;
		Dplus[585] = 12'b000000_000000;
		Dplus[586] = 12'b000000_000000;
		Dplus[587] = 12'b000000_000000;
		Dplus[588] = 12'b000000_000000;
		Dplus[589] = 12'b000000_000000;
		Dplus[590] = 12'b000000_000000;
		Dplus[591] = 12'b000000_000000;
		Dplus[592] = 12'b000000_000000;
		Dplus[593] = 12'b000000_000000;
		Dplus[594] = 12'b000000_000000;
		Dplus[595] = 12'b000000_000000;
		Dplus[596] = 12'b000000_000000;
		Dplus[597] = 12'b000000_000000;
		Dplus[598] = 12'b000000_000000;
		Dplus[599] = 12'b000000_000000;
		Dplus[600] = 12'b000000_000000;
		Dplus[601] = 12'b000000_000000;
		Dplus[602] = 12'b000000_000000;
		Dplus[603] = 12'b000000_000000;
		Dplus[604] = 12'b000000_000000;
		Dplus[605] = 12'b000000_000000;
		Dplus[606] = 12'b000000_000000;
		Dplus[607] = 12'b000000_000000;
		Dplus[608] = 12'b000000_000000;
		Dplus[609] = 12'b000000_000000;
		Dplus[610] = 12'b000000_000000;
		Dplus[611] = 12'b000000_000000;
		Dplus[612] = 12'b000000_000000;
		Dplus[613] = 12'b000000_000000;
		Dplus[614] = 12'b000000_000000;
		Dplus[615] = 12'b000000_000000;
		Dplus[616] = 12'b000000_000000;
		Dplus[617] = 12'b000000_000000;
		Dplus[618] = 12'b000000_000000;
		Dplus[619] = 12'b000000_000000;
		Dplus[620] = 12'b000000_000000;
		Dplus[621] = 12'b000000_000000;
		Dplus[622] = 12'b000000_000000;
		Dplus[623] = 12'b000000_000000;
		Dplus[624] = 12'b000000_000000;
		Dplus[625] = 12'b000000_000000;
		Dplus[626] = 12'b000000_000000;
		Dplus[627] = 12'b000000_000000;
		Dplus[628] = 12'b000000_000000;
		Dplus[629] = 12'b000000_000000;
		Dplus[630] = 12'b000000_000000;
		Dplus[631] = 12'b000000_000000;
		Dplus[632] = 12'b000000_000000;
		Dplus[633] = 12'b000000_000000;
		Dplus[634] = 12'b000000_000000;
		Dplus[635] = 12'b000000_000000;
		Dplus[636] = 12'b000000_000000;
		Dplus[637] = 12'b000000_000000;
		Dplus[638] = 12'b000000_000000;
		Dplus[639] = 12'b000000_000000;
		Dplus[640] = 12'b000000_000000;
		Dplus[641] = 12'b000000_000000;
		Dplus[642] = 12'b000000_000000;
		Dplus[643] = 12'b000000_000000;
		Dplus[644] = 12'b000000_000000;
		Dplus[645] = 12'b000000_000000;
		Dplus[646] = 12'b000000_000000;
		Dplus[647] = 12'b000000_000000;
		Dplus[648] = 12'b000000_000000;
		Dplus[649] = 12'b000000_000000;
		Dplus[650] = 12'b000000_000000;
		Dplus[651] = 12'b000000_000000;
		Dplus[652] = 12'b000000_000000;
		Dplus[653] = 12'b000000_000000;
		Dplus[654] = 12'b000000_000000;
		Dplus[655] = 12'b000000_000000;
		Dplus[656] = 12'b000000_000000;
		Dplus[657] = 12'b000000_000000;
		Dplus[658] = 12'b000000_000000;
		Dplus[659] = 12'b000000_000000;
		Dplus[660] = 12'b000000_000000;
		Dplus[661] = 12'b000000_000000;
		Dplus[662] = 12'b000000_000000;
		Dplus[663] = 12'b000000_000000;
		Dplus[664] = 12'b000000_000000;
		Dplus[665] = 12'b000000_000000;
		Dplus[666] = 12'b000000_000000;
		Dplus[667] = 12'b000000_000000;
		Dplus[668] = 12'b000000_000000;
		Dplus[669] = 12'b000000_000000;
		Dplus[670] = 12'b000000_000000;
		Dplus[671] = 12'b000000_000000;
		Dplus[672] = 12'b000000_000000;
		Dplus[673] = 12'b000000_000000;
		Dplus[674] = 12'b000000_000000;
		Dplus[675] = 12'b000000_000000;
		Dplus[676] = 12'b000000_000000;
		Dplus[677] = 12'b000000_000000;
		Dplus[678] = 12'b000000_000000;
		Dplus[679] = 12'b000000_000000;
		Dplus[680] = 12'b000000_000000;
		Dplus[681] = 12'b000000_000000;
		Dplus[682] = 12'b000000_000000;
		Dplus[683] = 12'b000000_000000;
		Dplus[684] = 12'b000000_000000;
		Dplus[685] = 12'b000000_000000;
		Dplus[686] = 12'b000000_000000;
		Dplus[687] = 12'b000000_000000;
		Dplus[688] = 12'b000000_000000;
		Dplus[689] = 12'b000000_000000;
		Dplus[690] = 12'b000000_000000;
		Dplus[691] = 12'b000000_000000;
		Dplus[692] = 12'b000000_000000;
		Dplus[693] = 12'b000000_000000;
		Dplus[694] = 12'b000000_000000;
		Dplus[695] = 12'b000000_000000;
		Dplus[696] = 12'b000000_000000;
		Dplus[697] = 12'b000000_000000;
		Dplus[698] = 12'b000000_000000;
		Dplus[699] = 12'b000000_000000;
		Dplus[700] = 12'b000000_000000;
		Dplus[701] = 12'b000000_000000;
		Dplus[702] = 12'b000000_000000;
		Dplus[703] = 12'b000000_000000;
		Dplus[704] = 12'b000000_000000;
		Dplus[705] = 12'b000000_000000;
		Dplus[706] = 12'b000000_000000;
		Dplus[707] = 12'b000000_000000;
		Dplus[708] = 12'b000000_000000;
		Dplus[709] = 12'b000000_000000;
		Dplus[710] = 12'b000000_000000;
		Dplus[711] = 12'b000000_000000;
		Dplus[712] = 12'b000000_000000;
		Dplus[713] = 12'b000000_000000;
		Dplus[714] = 12'b000000_000000;
		Dplus[715] = 12'b000000_000000;
		Dplus[716] = 12'b000000_000000;
		Dplus[717] = 12'b000000_000000;
		Dplus[718] = 12'b000000_000000;
		Dplus[719] = 12'b000000_000000;
		Dplus[720] = 12'b000000_000000;
		Dplus[721] = 12'b000000_000000;
		Dplus[722] = 12'b000000_000000;
		Dplus[723] = 12'b000000_000000;
		Dplus[724] = 12'b000000_000000;
		Dplus[725] = 12'b000000_000000;
		Dplus[726] = 12'b000000_000000;
		Dplus[727] = 12'b000000_000000;
		Dplus[728] = 12'b000000_000000;
		Dplus[729] = 12'b000000_000000;
		Dplus[730] = 12'b000000_000000;
		Dplus[731] = 12'b000000_000000;
		Dplus[732] = 12'b000000_000000;
		Dplus[733] = 12'b000000_000000;
		Dplus[734] = 12'b000000_000000;
		Dplus[735] = 12'b000000_000000;
		Dplus[736] = 12'b000000_000000;
		Dplus[737] = 12'b000000_000000;
		Dplus[738] = 12'b000000_000000;
		Dplus[739] = 12'b000000_000000;
		Dplus[740] = 12'b000000_000000;
		Dplus[741] = 12'b000000_000000;
		Dplus[742] = 12'b000000_000000;
		Dplus[743] = 12'b000000_000000;
		Dplus[744] = 12'b000000_000000;
		Dplus[745] = 12'b000000_000000;
		Dplus[746] = 12'b000000_000000;
		Dplus[747] = 12'b000000_000000;
		Dplus[748] = 12'b000000_000000;
		Dplus[749] = 12'b000000_000000;
		Dplus[750] = 12'b000000_000000;
		Dplus[751] = 12'b000000_000000;
		Dplus[752] = 12'b000000_000000;
		Dplus[753] = 12'b000000_000000;
		Dplus[754] = 12'b000000_000000;
		Dplus[755] = 12'b000000_000000;
		Dplus[756] = 12'b000000_000000;
		Dplus[757] = 12'b000000_000000;
		Dplus[758] = 12'b000000_000000;
		Dplus[759] = 12'b000000_000000;
		Dplus[760] = 12'b000000_000000;
		Dplus[761] = 12'b000000_000000;
		Dplus[762] = 12'b000000_000000;
		Dplus[763] = 12'b000000_000000;
		Dplus[764] = 12'b000000_000000;
		Dplus[765] = 12'b000000_000000;
		Dplus[766] = 12'b000000_000000;
		Dplus[767] = 12'b000000_000000;
		Dplus[768] = 12'b000000_000000;
		Dplus[769] = 12'b000000_000000;
		Dplus[770] = 12'b000000_000000;
		Dplus[771] = 12'b000000_000000;
		Dplus[772] = 12'b000000_000000;
		Dplus[773] = 12'b000000_000000;
		Dplus[774] = 12'b000000_000000;
		Dplus[775] = 12'b000000_000000;
		Dplus[776] = 12'b000000_000000;
		Dplus[777] = 12'b000000_000000;
		Dplus[778] = 12'b000000_000000;
		Dplus[779] = 12'b000000_000000;
		Dplus[780] = 12'b000000_000000;
		Dplus[781] = 12'b000000_000000;
		Dplus[782] = 12'b000000_000000;
		Dplus[783] = 12'b000000_000000;
		Dplus[784] = 12'b000000_000000;
		Dplus[785] = 12'b000000_000000;
		Dplus[786] = 12'b000000_000000;
		Dplus[787] = 12'b000000_000000;
		Dplus[788] = 12'b000000_000000;
		Dplus[789] = 12'b000000_000000;
		Dplus[790] = 12'b000000_000000;
		Dplus[791] = 12'b000000_000000;
		Dplus[792] = 12'b000000_000000;
		Dplus[793] = 12'b000000_000000;
		Dplus[794] = 12'b000000_000000;
		Dplus[795] = 12'b000000_000000;
		Dplus[796] = 12'b000000_000000;
		Dplus[797] = 12'b000000_000000;
		Dplus[798] = 12'b000000_000000;
		Dplus[799] = 12'b000000_000000;
		Dplus[800] = 12'b000000_000000;
		Dplus[801] = 12'b000000_000000;
		Dplus[802] = 12'b000000_000000;
		Dplus[803] = 12'b000000_000000;
		Dplus[804] = 12'b000000_000000;
		Dplus[805] = 12'b000000_000000;
		Dplus[806] = 12'b000000_000000;
		Dplus[807] = 12'b000000_000000;
		Dplus[808] = 12'b000000_000000;
		Dplus[809] = 12'b000000_000000;
		Dplus[810] = 12'b000000_000000;
		Dplus[811] = 12'b000000_000000;
		Dplus[812] = 12'b000000_000000;
		Dplus[813] = 12'b000000_000000;
		Dplus[814] = 12'b000000_000000;
		Dplus[815] = 12'b000000_000000;
		Dplus[816] = 12'b000000_000000;
		Dplus[817] = 12'b000000_000000;
		Dplus[818] = 12'b000000_000000;
		Dplus[819] = 12'b000000_000000;
		Dplus[820] = 12'b000000_000000;
		Dplus[821] = 12'b000000_000000;
		Dplus[822] = 12'b000000_000000;
		Dplus[823] = 12'b000000_000000;
		Dplus[824] = 12'b000000_000000;
		Dplus[825] = 12'b000000_000000;
		Dplus[826] = 12'b000000_000000;
		Dplus[827] = 12'b000000_000000;
		Dplus[828] = 12'b000000_000000;
		Dplus[829] = 12'b000000_000000;
		Dplus[830] = 12'b000000_000000;
		Dplus[831] = 12'b000000_000000;
		Dplus[832] = 12'b000000_000000;
		Dplus[833] = 12'b000000_000000;
		Dplus[834] = 12'b000000_000000;
		Dplus[835] = 12'b000000_000000;
		Dplus[836] = 12'b000000_000000;
		Dplus[837] = 12'b000000_000000;
		Dplus[838] = 12'b000000_000000;
		Dplus[839] = 12'b000000_000000;
		Dplus[840] = 12'b000000_000000;
		Dplus[841] = 12'b000000_000000;
		Dplus[842] = 12'b000000_000000;
		Dplus[843] = 12'b000000_000000;
		Dplus[844] = 12'b000000_000000;
		Dplus[845] = 12'b000000_000000;
		Dplus[846] = 12'b000000_000000;
		Dplus[847] = 12'b000000_000000;
		Dplus[848] = 12'b000000_000000;
		Dplus[849] = 12'b000000_000000;
		Dplus[850] = 12'b000000_000000;
		Dplus[851] = 12'b000000_000000;
		Dplus[852] = 12'b000000_000000;
		Dplus[853] = 12'b000000_000000;
		Dplus[854] = 12'b000000_000000;
		Dplus[855] = 12'b000000_000000;
		Dplus[856] = 12'b000000_000000;
		Dplus[857] = 12'b000000_000000;
		Dplus[858] = 12'b000000_000000;
		Dplus[859] = 12'b000000_000000;
		Dplus[860] = 12'b000000_000000;
		Dplus[861] = 12'b000000_000000;
		Dplus[862] = 12'b000000_000000;
		Dplus[863] = 12'b000000_000000;
		Dplus[864] = 12'b000000_000000;
		Dplus[865] = 12'b000000_000000;
		Dplus[866] = 12'b000000_000000;
		Dplus[867] = 12'b000000_000000;
		Dplus[868] = 12'b000000_000000;
		Dplus[869] = 12'b000000_000000;
		Dplus[870] = 12'b000000_000000;
		Dplus[871] = 12'b000000_000000;
		Dplus[872] = 12'b000000_000000;
		Dplus[873] = 12'b000000_000000;
		Dplus[874] = 12'b000000_000000;
		Dplus[875] = 12'b000000_000000;
		Dplus[876] = 12'b000000_000000;
		Dplus[877] = 12'b000000_000000;
		Dplus[878] = 12'b000000_000000;
		Dplus[879] = 12'b000000_000000;
		Dplus[880] = 12'b000000_000000;
		Dplus[881] = 12'b000000_000000;
		Dplus[882] = 12'b000000_000000;
		Dplus[883] = 12'b000000_000000;
		Dplus[884] = 12'b000000_000000;
		Dplus[885] = 12'b000000_000000;
		Dplus[886] = 12'b000000_000000;
		Dplus[887] = 12'b000000_000000;
		Dplus[888] = 12'b000000_000000;
		Dplus[889] = 12'b000000_000000;
		Dplus[890] = 12'b000000_000000;
		Dplus[891] = 12'b000000_000000;
		Dplus[892] = 12'b000000_000000;
		Dplus[893] = 12'b000000_000000;
		Dplus[894] = 12'b000000_000000;
		Dplus[895] = 12'b000000_000000;
		Dplus[896] = 12'b000000_000000;
		Dplus[897] = 12'b000000_000000;
		Dplus[898] = 12'b000000_000000;
		Dplus[899] = 12'b000000_000000;
		Dplus[900] = 12'b000000_000000;
		Dplus[901] = 12'b000000_000000;
		Dplus[902] = 12'b000000_000000;
		Dplus[903] = 12'b000000_000000;
		Dplus[904] = 12'b000000_000000;
		Dplus[905] = 12'b000000_000000;
		Dplus[906] = 12'b000000_000000;
		Dplus[907] = 12'b000000_000000;
		Dplus[908] = 12'b000000_000000;
		Dplus[909] = 12'b000000_000000;
		Dplus[910] = 12'b000000_000000;
		Dplus[911] = 12'b000000_000000;
		Dplus[912] = 12'b000000_000000;
		Dplus[913] = 12'b000000_000000;
		Dplus[914] = 12'b000000_000000;
		Dplus[915] = 12'b000000_000000;
		Dplus[916] = 12'b000000_000000;
		Dplus[917] = 12'b000000_000000;
		Dplus[918] = 12'b000000_000000;
		Dplus[919] = 12'b000000_000000;
		Dplus[920] = 12'b000000_000000;
		Dplus[921] = 12'b000000_000000;
		Dplus[922] = 12'b000000_000000;
		Dplus[923] = 12'b000000_000000;
		Dplus[924] = 12'b000000_000000;
		Dplus[925] = 12'b000000_000000;
		Dplus[926] = 12'b000000_000000;
		Dplus[927] = 12'b000000_000000;
		Dplus[928] = 12'b000000_000000;
		Dplus[929] = 12'b000000_000000;
		Dplus[930] = 12'b000000_000000;
		Dplus[931] = 12'b000000_000000;
		Dplus[932] = 12'b000000_000000;
		Dplus[933] = 12'b000000_000000;
		Dplus[934] = 12'b000000_000000;
		Dplus[935] = 12'b000000_000000;
		Dplus[936] = 12'b000000_000000;
		Dplus[937] = 12'b000000_000000;
		Dplus[938] = 12'b000000_000000;
		Dplus[939] = 12'b000000_000000;
		Dplus[940] = 12'b000000_000000;
		Dplus[941] = 12'b000000_000000;
		Dplus[942] = 12'b000000_000000;
		Dplus[943] = 12'b000000_000000;
		Dplus[944] = 12'b000000_000000;
		Dplus[945] = 12'b000000_000000;
		Dplus[946] = 12'b000000_000000;
		Dplus[947] = 12'b000000_000000;
		Dplus[948] = 12'b000000_000000;
		Dplus[949] = 12'b000000_000000;
		Dplus[950] = 12'b000000_000000;
		Dplus[951] = 12'b000000_000000;
		Dplus[952] = 12'b000000_000000;
		Dplus[953] = 12'b000000_000000;
		Dplus[954] = 12'b000000_000000;
		Dplus[955] = 12'b000000_000000;
		Dplus[956] = 12'b000000_000000;
		Dplus[957] = 12'b000000_000000;
		Dplus[958] = 12'b000000_000000;
		Dplus[959] = 12'b000000_000000;
		Dplus[960] = 12'b000000_000000;
		Dplus[961] = 12'b000000_000000;
		Dplus[962] = 12'b000000_000000;
		Dplus[963] = 12'b000000_000000;
		Dplus[964] = 12'b000000_000000;
		Dplus[965] = 12'b000000_000000;
		Dplus[966] = 12'b000000_000000;
		Dplus[967] = 12'b000000_000000;
		Dplus[968] = 12'b000000_000000;
		Dplus[969] = 12'b000000_000000;
		Dplus[970] = 12'b000000_000000;
		Dplus[971] = 12'b000000_000000;
		Dplus[972] = 12'b000000_000000;
		Dplus[973] = 12'b000000_000000;
		Dplus[974] = 12'b000000_000000;
		Dplus[975] = 12'b000000_000000;
		Dplus[976] = 12'b000000_000000;
		Dplus[977] = 12'b000000_000000;
		Dplus[978] = 12'b000000_000000;
		Dplus[979] = 12'b000000_000000;
		Dplus[980] = 12'b000000_000000;
		Dplus[981] = 12'b000000_000000;
		Dplus[982] = 12'b000000_000000;
		Dplus[983] = 12'b000000_000000;
		Dplus[984] = 12'b000000_000000;
		Dplus[985] = 12'b000000_000000;
		Dplus[986] = 12'b000000_000000;
		Dplus[987] = 12'b000000_000000;
		Dplus[988] = 12'b000000_000000;
		Dplus[989] = 12'b000000_000000;
		Dplus[990] = 12'b000000_000000;
		Dplus[991] = 12'b000000_000000;
		Dplus[992] = 12'b000000_000000;
		Dplus[993] = 12'b000000_000000;
		Dplus[994] = 12'b000000_000000;
		Dplus[995] = 12'b000000_000000;
		Dplus[996] = 12'b000000_000000;
		Dplus[997] = 12'b000000_000000;
		Dplus[998] = 12'b000000_000000;
		Dplus[999] = 12'b000000_000000;
		Dplus[1000] = 12'b000000_000000;
		Dplus[1001] = 12'b000000_000000;
		Dplus[1002] = 12'b000000_000000;
		Dplus[1003] = 12'b000000_000000;
		Dplus[1004] = 12'b000000_000000;
		Dplus[1005] = 12'b000000_000000;
		Dplus[1006] = 12'b000000_000000;
		Dplus[1007] = 12'b000000_000000;
		Dplus[1008] = 12'b000000_000000;
		Dplus[1009] = 12'b000000_000000;
		Dplus[1010] = 12'b000000_000000;
		Dplus[1011] = 12'b000000_000000;
		Dplus[1012] = 12'b000000_000000;
		Dplus[1013] = 12'b000000_000000;
		Dplus[1014] = 12'b000000_000000;
		Dplus[1015] = 12'b000000_000000;
		Dplus[1016] = 12'b000000_000000;
		Dplus[1017] = 12'b000000_000000;
		Dplus[1018] = 12'b000000_000000;
		Dplus[1019] = 12'b000000_000000;
		Dplus[1020] = 12'b000000_000000;
		Dplus[1021] = 12'b000000_000000;
		Dplus[1022] = 12'b000000_000000;
		Dplus[1023] = 12'b000000_000000;
		Dplus[1024] = 12'b000000_000000;
		Dplus[1025] = 12'b000000_000000;
		Dplus[1026] = 12'b000000_000000;
		Dplus[1027] = 12'b000000_000000;
		Dplus[1028] = 12'b000000_000000;
		Dplus[1029] = 12'b000000_000000;
		Dplus[1030] = 12'b000000_000000;
		Dplus[1031] = 12'b000000_000000;
		Dplus[1032] = 12'b000000_000000;
		Dplus[1033] = 12'b000000_000000;
		Dplus[1034] = 12'b000000_000000;
		Dplus[1035] = 12'b000000_000000;
		Dplus[1036] = 12'b000000_000000;
		Dplus[1037] = 12'b000000_000000;
		Dplus[1038] = 12'b000000_000000;
		Dplus[1039] = 12'b000000_000000;
		Dplus[1040] = 12'b000000_000000;
		Dplus[1041] = 12'b000000_000000;
		Dplus[1042] = 12'b000000_000000;
		Dplus[1043] = 12'b000000_000000;
		Dplus[1044] = 12'b000000_000000;
		Dplus[1045] = 12'b000000_000000;
		Dplus[1046] = 12'b000000_000000;
		Dplus[1047] = 12'b000000_000000;
		Dplus[1048] = 12'b000000_000000;
		Dplus[1049] = 12'b000000_000000;
		Dplus[1050] = 12'b000000_000000;
		Dplus[1051] = 12'b000000_000000;
		Dplus[1052] = 12'b000000_000000;
		Dplus[1053] = 12'b000000_000000;
		Dplus[1054] = 12'b000000_000000;
		Dplus[1055] = 12'b000000_000000;
		Dplus[1056] = 12'b000000_000000;
		Dplus[1057] = 12'b000000_000000;
		Dplus[1058] = 12'b000000_000000;
		Dplus[1059] = 12'b000000_000000;
		Dplus[1060] = 12'b000000_000000;
		Dplus[1061] = 12'b000000_000000;
		Dplus[1062] = 12'b000000_000000;
		Dplus[1063] = 12'b000000_000000;
		Dplus[1064] = 12'b000000_000000;
		Dplus[1065] = 12'b000000_000000;
		Dplus[1066] = 12'b000000_000000;
		Dplus[1067] = 12'b000000_000000;
		Dplus[1068] = 12'b000000_000000;
		Dplus[1069] = 12'b000000_000000;
		Dplus[1070] = 12'b000000_000000;
		Dplus[1071] = 12'b000000_000000;
		Dplus[1072] = 12'b000000_000000;
		Dplus[1073] = 12'b000000_000000;
		Dplus[1074] = 12'b000000_000000;
		Dplus[1075] = 12'b000000_000000;
		Dplus[1076] = 12'b000000_000000;
		Dplus[1077] = 12'b000000_000000;
		Dplus[1078] = 12'b000000_000000;
		Dplus[1079] = 12'b000000_000000;
		Dplus[1080] = 12'b000000_000000;
		Dplus[1081] = 12'b000000_000000;
		Dplus[1082] = 12'b000000_000000;
		Dplus[1083] = 12'b000000_000000;
		Dplus[1084] = 12'b000000_000000;
		Dplus[1085] = 12'b000000_000000;
		Dplus[1086] = 12'b000000_000000;
		Dplus[1087] = 12'b000000_000000;
		Dplus[1088] = 12'b000000_000000;
		Dplus[1089] = 12'b000000_000000;
		Dplus[1090] = 12'b000000_000000;
		Dplus[1091] = 12'b000000_000000;
		Dplus[1092] = 12'b000000_000000;
		Dplus[1093] = 12'b000000_000000;
		Dplus[1094] = 12'b000000_000000;
		Dplus[1095] = 12'b000000_000000;
		Dplus[1096] = 12'b000000_000000;
		Dplus[1097] = 12'b000000_000000;
		Dplus[1098] = 12'b000000_000000;
		Dplus[1099] = 12'b000000_000000;
		Dplus[1100] = 12'b000000_000000;
		Dplus[1101] = 12'b000000_000000;
		Dplus[1102] = 12'b000000_000000;
		Dplus[1103] = 12'b000000_000000;
		Dplus[1104] = 12'b000000_000000;
		Dplus[1105] = 12'b000000_000000;
		Dplus[1106] = 12'b000000_000000;
		Dplus[1107] = 12'b000000_000000;
		Dplus[1108] = 12'b000000_000000;
		Dplus[1109] = 12'b000000_000000;
		Dplus[1110] = 12'b000000_000000;
		Dplus[1111] = 12'b000000_000000;
		Dplus[1112] = 12'b000000_000000;
		Dplus[1113] = 12'b000000_000000;
		Dplus[1114] = 12'b000000_000000;
		Dplus[1115] = 12'b000000_000000;
		Dplus[1116] = 12'b000000_000000;
		Dplus[1117] = 12'b000000_000000;
		Dplus[1118] = 12'b000000_000000;
		Dplus[1119] = 12'b000000_000000;
		Dplus[1120] = 12'b000000_000000;
		Dplus[1121] = 12'b000000_000000;
		Dplus[1122] = 12'b000000_000000;
		Dplus[1123] = 12'b000000_000000;
		Dplus[1124] = 12'b000000_000000;
		Dplus[1125] = 12'b000000_000000;
		Dplus[1126] = 12'b000000_000000;
		Dplus[1127] = 12'b000000_000000;
		Dplus[1128] = 12'b000000_000000;
		Dplus[1129] = 12'b000000_000000;
		Dplus[1130] = 12'b000000_000000;
		Dplus[1131] = 12'b000000_000000;
		Dplus[1132] = 12'b000000_000000;
		Dplus[1133] = 12'b000000_000000;
		Dplus[1134] = 12'b000000_000000;
		Dplus[1135] = 12'b000000_000000;
		Dplus[1136] = 12'b000000_000000;
		Dplus[1137] = 12'b000000_000000;
		Dplus[1138] = 12'b000000_000000;
		Dplus[1139] = 12'b000000_000000;
		Dplus[1140] = 12'b000000_000000;
		Dplus[1141] = 12'b000000_000000;
		Dplus[1142] = 12'b000000_000000;
		Dplus[1143] = 12'b000000_000000;
		Dplus[1144] = 12'b000000_000000;
		Dplus[1145] = 12'b000000_000000;
		Dplus[1146] = 12'b000000_000000;
		Dplus[1147] = 12'b000000_000000;
		Dplus[1148] = 12'b000000_000000;
		Dplus[1149] = 12'b000000_000000;
		Dplus[1150] = 12'b000000_000000;
		Dplus[1151] = 12'b000000_000000;
		Dplus[1152] = 12'b000000_000000;
		Dplus[1153] = 12'b000000_000000;
		Dplus[1154] = 12'b000000_000000;
		Dplus[1155] = 12'b000000_000000;
		Dplus[1156] = 12'b000000_000000;
		Dplus[1157] = 12'b000000_000000;
		Dplus[1158] = 12'b000000_000000;
		Dplus[1159] = 12'b000000_000000;
		Dplus[1160] = 12'b000000_000000;
		Dplus[1161] = 12'b000000_000000;
		Dplus[1162] = 12'b000000_000000;
		Dplus[1163] = 12'b000000_000000;
		Dplus[1164] = 12'b000000_000000;
		Dplus[1165] = 12'b000000_000000;
		Dplus[1166] = 12'b000000_000000;
		Dplus[1167] = 12'b000000_000000;
		Dplus[1168] = 12'b000000_000000;
		Dplus[1169] = 12'b000000_000000;
		Dplus[1170] = 12'b000000_000000;
		Dplus[1171] = 12'b000000_000000;
		Dplus[1172] = 12'b000000_000000;
		Dplus[1173] = 12'b000000_000000;
		Dplus[1174] = 12'b000000_000000;
		Dplus[1175] = 12'b000000_000000;
		Dplus[1176] = 12'b000000_000000;
		Dplus[1177] = 12'b000000_000000;
		Dplus[1178] = 12'b000000_000000;
		Dplus[1179] = 12'b000000_000000;
		Dplus[1180] = 12'b000000_000000;
		Dplus[1181] = 12'b000000_000000;
		Dplus[1182] = 12'b000000_000000;
		Dplus[1183] = 12'b000000_000000;
		Dplus[1184] = 12'b000000_000000;
		Dplus[1185] = 12'b000000_000000;
		Dplus[1186] = 12'b000000_000000;
		Dplus[1187] = 12'b000000_000000;
		Dplus[1188] = 12'b000000_000000;
		Dplus[1189] = 12'b000000_000000;
		Dplus[1190] = 12'b000000_000000;
		Dplus[1191] = 12'b000000_000000;
		Dplus[1192] = 12'b000000_000000;
		Dplus[1193] = 12'b000000_000000;
		Dplus[1194] = 12'b000000_000000;
		Dplus[1195] = 12'b000000_000000;
		Dplus[1196] = 12'b000000_000000;
		Dplus[1197] = 12'b000000_000000;
		Dplus[1198] = 12'b000000_000000;
		Dplus[1199] = 12'b000000_000000;
		Dplus[1200] = 12'b000000_000000;
		Dplus[1201] = 12'b000000_000000;
		Dplus[1202] = 12'b000000_000000;
		Dplus[1203] = 12'b000000_000000;
		Dplus[1204] = 12'b000000_000000;
		Dplus[1205] = 12'b000000_000000;
		Dplus[1206] = 12'b000000_000000;
		Dplus[1207] = 12'b000000_000000;
		Dplus[1208] = 12'b000000_000000;
		Dplus[1209] = 12'b000000_000000;
		Dplus[1210] = 12'b000000_000000;
		Dplus[1211] = 12'b000000_000000;
		Dplus[1212] = 12'b000000_000000;
		Dplus[1213] = 12'b000000_000000;
		Dplus[1214] = 12'b000000_000000;
		Dplus[1215] = 12'b000000_000000;
		Dplus[1216] = 12'b000000_000000;
		Dplus[1217] = 12'b000000_000000;
		Dplus[1218] = 12'b000000_000000;
		Dplus[1219] = 12'b000000_000000;
		Dplus[1220] = 12'b000000_000000;
		Dplus[1221] = 12'b000000_000000;
		Dplus[1222] = 12'b000000_000000;
		Dplus[1223] = 12'b000000_000000;
		Dplus[1224] = 12'b000000_000000;
		Dplus[1225] = 12'b000000_000000;
		Dplus[1226] = 12'b000000_000000;
		Dplus[1227] = 12'b000000_000000;
		Dplus[1228] = 12'b000000_000000;
		Dplus[1229] = 12'b000000_000000;
		Dplus[1230] = 12'b000000_000000;
		Dplus[1231] = 12'b000000_000000;
		Dplus[1232] = 12'b000000_000000;
		Dplus[1233] = 12'b000000_000000;
		Dplus[1234] = 12'b000000_000000;
		Dplus[1235] = 12'b000000_000000;
		Dplus[1236] = 12'b000000_000000;
		Dplus[1237] = 12'b000000_000000;
		Dplus[1238] = 12'b000000_000000;
		Dplus[1239] = 12'b000000_000000;
		Dplus[1240] = 12'b000000_000000;
		Dplus[1241] = 12'b000000_000000;
		Dplus[1242] = 12'b000000_000000;
		Dplus[1243] = 12'b000000_000000;
		Dplus[1244] = 12'b000000_000000;
		Dplus[1245] = 12'b000000_000000;
		Dplus[1246] = 12'b000000_000000;
		Dplus[1247] = 12'b000000_000000;
		Dplus[1248] = 12'b000000_000000;
		Dplus[1249] = 12'b000000_000000;
		Dplus[1250] = 12'b000000_000000;
		Dplus[1251] = 12'b000000_000000;
		Dplus[1252] = 12'b000000_000000;
		Dplus[1253] = 12'b000000_000000;
		Dplus[1254] = 12'b000000_000000;
		Dplus[1255] = 12'b000000_000000;
		Dplus[1256] = 12'b000000_000000;
		Dplus[1257] = 12'b000000_000000;
		Dplus[1258] = 12'b000000_000000;
		Dplus[1259] = 12'b000000_000000;
		Dplus[1260] = 12'b000000_000000;
		Dplus[1261] = 12'b000000_000000;
		Dplus[1262] = 12'b000000_000000;
		Dplus[1263] = 12'b000000_000000;
		Dplus[1264] = 12'b000000_000000;
		Dplus[1265] = 12'b000000_000000;
		Dplus[1266] = 12'b000000_000000;
		Dplus[1267] = 12'b000000_000000;
		Dplus[1268] = 12'b000000_000000;
		Dplus[1269] = 12'b000000_000000;
		Dplus[1270] = 12'b000000_000000;
		Dplus[1271] = 12'b000000_000000;
		Dplus[1272] = 12'b000000_000000;
		Dplus[1273] = 12'b000000_000000;
		Dplus[1274] = 12'b000000_000000;
		Dplus[1275] = 12'b000000_000000;
		Dplus[1276] = 12'b000000_000000;
		Dplus[1277] = 12'b000000_000000;
		Dplus[1278] = 12'b000000_000000;
		Dplus[1279] = 12'b000000_000000;
		Dplus[1280] = 12'b000000_000000;
		Dplus[1281] = 12'b000000_000000;
		Dplus[1282] = 12'b000000_000000;
		Dplus[1283] = 12'b000000_000000;
		Dplus[1284] = 12'b000000_000000;
		Dplus[1285] = 12'b000000_000000;
		Dplus[1286] = 12'b000000_000000;
		Dplus[1287] = 12'b000000_000000;
		Dplus[1288] = 12'b000000_000000;
		Dplus[1289] = 12'b000000_000000;
		Dplus[1290] = 12'b000000_000000;
		Dplus[1291] = 12'b000000_000000;
		Dplus[1292] = 12'b000000_000000;
		Dplus[1293] = 12'b000000_000000;
		Dplus[1294] = 12'b000000_000000;
		Dplus[1295] = 12'b000000_000000;
		Dplus[1296] = 12'b000000_000000;
		Dplus[1297] = 12'b000000_000000;
		Dplus[1298] = 12'b000000_000000;
		Dplus[1299] = 12'b000000_000000;
		Dplus[1300] = 12'b000000_000000;
		Dplus[1301] = 12'b000000_000000;
		Dplus[1302] = 12'b000000_000000;
		Dplus[1303] = 12'b000000_000000;
		Dplus[1304] = 12'b000000_000000;
		Dplus[1305] = 12'b000000_000000;
		Dplus[1306] = 12'b000000_000000;
		Dplus[1307] = 12'b000000_000000;
		Dplus[1308] = 12'b000000_000000;
		Dplus[1309] = 12'b000000_000000;
		Dplus[1310] = 12'b000000_000000;
		Dplus[1311] = 12'b000000_000000;
		Dplus[1312] = 12'b000000_000000;
		Dplus[1313] = 12'b000000_000000;
		Dplus[1314] = 12'b000000_000000;
		Dplus[1315] = 12'b000000_000000;
		Dplus[1316] = 12'b000000_000000;
		Dplus[1317] = 12'b000000_000000;
		Dplus[1318] = 12'b000000_000000;
		Dplus[1319] = 12'b000000_000000;
		Dplus[1320] = 12'b000000_000000;
		Dplus[1321] = 12'b000000_000000;
		Dplus[1322] = 12'b000000_000000;
		Dplus[1323] = 12'b000000_000000;
		Dplus[1324] = 12'b000000_000000;
		Dplus[1325] = 12'b000000_000000;
		Dplus[1326] = 12'b000000_000000;
		Dplus[1327] = 12'b000000_000000;
		Dplus[1328] = 12'b000000_000000;
		Dplus[1329] = 12'b000000_000000;
		Dplus[1330] = 12'b000000_000000;
		Dplus[1331] = 12'b000000_000000;
		Dplus[1332] = 12'b000000_000000;
		Dplus[1333] = 12'b000000_000000;
		Dplus[1334] = 12'b000000_000000;
		Dplus[1335] = 12'b000000_000000;
		Dplus[1336] = 12'b000000_000000;
		Dplus[1337] = 12'b000000_000000;
		Dplus[1338] = 12'b000000_000000;
		Dplus[1339] = 12'b000000_000000;
		Dplus[1340] = 12'b000000_000000;
		Dplus[1341] = 12'b000000_000000;
		Dplus[1342] = 12'b000000_000000;
		Dplus[1343] = 12'b000000_000000;
		Dplus[1344] = 12'b000000_000000;
		Dplus[1345] = 12'b000000_000000;
		Dplus[1346] = 12'b000000_000000;
		Dplus[1347] = 12'b000000_000000;
		Dplus[1348] = 12'b000000_000000;
		Dplus[1349] = 12'b000000_000000;
		Dplus[1350] = 12'b000000_000000;
		Dplus[1351] = 12'b000000_000000;
		Dplus[1352] = 12'b000000_000000;
		Dplus[1353] = 12'b000000_000000;
		Dplus[1354] = 12'b000000_000000;
		Dplus[1355] = 12'b000000_000000;
		Dplus[1356] = 12'b000000_000000;
		Dplus[1357] = 12'b000000_000000;
		Dplus[1358] = 12'b000000_000000;
		Dplus[1359] = 12'b000000_000000;
		Dplus[1360] = 12'b000000_000000;
		Dplus[1361] = 12'b000000_000000;
		Dplus[1362] = 12'b000000_000000;
		Dplus[1363] = 12'b000000_000000;
		Dplus[1364] = 12'b000000_000000;
		Dplus[1365] = 12'b000000_000000;
		Dplus[1366] = 12'b000000_000000;
		Dplus[1367] = 12'b000000_000000;
		Dplus[1368] = 12'b000000_000000;
		Dplus[1369] = 12'b000000_000000;
		Dplus[1370] = 12'b000000_000000;
		Dplus[1371] = 12'b000000_000000;
		Dplus[1372] = 12'b000000_000000;
		Dplus[1373] = 12'b000000_000000;
		Dplus[1374] = 12'b000000_000000;
		Dplus[1375] = 12'b000000_000000;
		Dplus[1376] = 12'b000000_000000;
		Dplus[1377] = 12'b000000_000000;
		Dplus[1378] = 12'b000000_000000;
		Dplus[1379] = 12'b000000_000000;
		Dplus[1380] = 12'b000000_000000;
		Dplus[1381] = 12'b000000_000000;
		Dplus[1382] = 12'b000000_000000;
		Dplus[1383] = 12'b000000_000000;
		Dplus[1384] = 12'b000000_000000;
		Dplus[1385] = 12'b000000_000000;
		Dplus[1386] = 12'b000000_000000;
		Dplus[1387] = 12'b000000_000000;
		Dplus[1388] = 12'b000000_000000;
		Dplus[1389] = 12'b000000_000000;
		Dplus[1390] = 12'b000000_000000;
		Dplus[1391] = 12'b000000_000000;
		Dplus[1392] = 12'b000000_000000;
		Dplus[1393] = 12'b000000_000000;
		Dplus[1394] = 12'b000000_000000;
		Dplus[1395] = 12'b000000_000000;
		Dplus[1396] = 12'b000000_000000;
		Dplus[1397] = 12'b000000_000000;
		Dplus[1398] = 12'b000000_000000;
		Dplus[1399] = 12'b000000_000000;
		Dplus[1400] = 12'b000000_000000;
		Dplus[1401] = 12'b000000_000000;
		Dplus[1402] = 12'b000000_000000;
		Dplus[1403] = 12'b000000_000000;
		Dplus[1404] = 12'b000000_000000;
		Dplus[1405] = 12'b000000_000000;
		Dplus[1406] = 12'b000000_000000;
		Dplus[1407] = 12'b000000_000000;
		Dplus[1408] = 12'b000000_000000;
		Dplus[1409] = 12'b000000_000000;
		Dplus[1410] = 12'b000000_000000;
		Dplus[1411] = 12'b000000_000000;
		Dplus[1412] = 12'b000000_000000;
		Dplus[1413] = 12'b000000_000000;
		Dplus[1414] = 12'b000000_000000;
		Dplus[1415] = 12'b000000_000000;
		Dplus[1416] = 12'b000000_000000;
		Dplus[1417] = 12'b000000_000000;
		Dplus[1418] = 12'b000000_000000;
		Dplus[1419] = 12'b000000_000000;
		Dplus[1420] = 12'b000000_000000;
		Dplus[1421] = 12'b000000_000000;
		Dplus[1422] = 12'b000000_000000;
		Dplus[1423] = 12'b000000_000000;
		Dplus[1424] = 12'b000000_000000;
		Dplus[1425] = 12'b000000_000000;
		Dplus[1426] = 12'b000000_000000;
		Dplus[1427] = 12'b000000_000000;
		Dplus[1428] = 12'b000000_000000;
		Dplus[1429] = 12'b000000_000000;
		Dplus[1430] = 12'b000000_000000;
		Dplus[1431] = 12'b000000_000000;
		Dplus[1432] = 12'b000000_000000;
		Dplus[1433] = 12'b000000_000000;
		Dplus[1434] = 12'b000000_000000;
		Dplus[1435] = 12'b000000_000000;
		Dplus[1436] = 12'b000000_000000;
		Dplus[1437] = 12'b000000_000000;
		Dplus[1438] = 12'b000000_000000;
		Dplus[1439] = 12'b000000_000000;
		Dplus[1440] = 12'b000000_000000;
		Dplus[1441] = 12'b000000_000000;
		Dplus[1442] = 12'b000000_000000;
		Dplus[1443] = 12'b000000_000000;
		Dplus[1444] = 12'b000000_000000;
		Dplus[1445] = 12'b000000_000000;
		Dplus[1446] = 12'b000000_000000;
		Dplus[1447] = 12'b000000_000000;
		Dplus[1448] = 12'b000000_000000;
		Dplus[1449] = 12'b000000_000000;
		Dplus[1450] = 12'b000000_000000;
		Dplus[1451] = 12'b000000_000000;
		Dplus[1452] = 12'b000000_000000;
		Dplus[1453] = 12'b000000_000000;
		Dplus[1454] = 12'b000000_000000;
		Dplus[1455] = 12'b000000_000000;
		Dplus[1456] = 12'b000000_000000;
		Dplus[1457] = 12'b000000_000000;
		Dplus[1458] = 12'b000000_000000;
		Dplus[1459] = 12'b000000_000000;
		Dplus[1460] = 12'b000000_000000;
		Dplus[1461] = 12'b000000_000000;
		Dplus[1462] = 12'b000000_000000;
		Dplus[1463] = 12'b000000_000000;
		Dplus[1464] = 12'b000000_000000;
		Dplus[1465] = 12'b000000_000000;
		Dplus[1466] = 12'b000000_000000;
		Dplus[1467] = 12'b000000_000000;
		Dplus[1468] = 12'b000000_000000;
		Dplus[1469] = 12'b000000_000000;
		Dplus[1470] = 12'b000000_000000;
		Dplus[1471] = 12'b000000_000000;
		Dplus[1472] = 12'b000000_000000;
		Dplus[1473] = 12'b000000_000000;
		Dplus[1474] = 12'b000000_000000;
		Dplus[1475] = 12'b000000_000000;
		Dplus[1476] = 12'b000000_000000;
		Dplus[1477] = 12'b000000_000000;
		Dplus[1478] = 12'b000000_000000;
		Dplus[1479] = 12'b000000_000000;
		Dplus[1480] = 12'b000000_000000;
		Dplus[1481] = 12'b000000_000000;
		Dplus[1482] = 12'b000000_000000;
		Dplus[1483] = 12'b000000_000000;
		Dplus[1484] = 12'b000000_000000;
		Dplus[1485] = 12'b000000_000000;
		Dplus[1486] = 12'b000000_000000;
		Dplus[1487] = 12'b000000_000000;
		Dplus[1488] = 12'b000000_000000;
		Dplus[1489] = 12'b000000_000000;
		Dplus[1490] = 12'b000000_000000;
		Dplus[1491] = 12'b000000_000000;
		Dplus[1492] = 12'b000000_000000;
		Dplus[1493] = 12'b000000_000000;
		Dplus[1494] = 12'b000000_000000;
		Dplus[1495] = 12'b000000_000000;
		Dplus[1496] = 12'b000000_000000;
		Dplus[1497] = 12'b000000_000000;
		Dplus[1498] = 12'b000000_000000;
		Dplus[1499] = 12'b000000_000000;
		Dplus[1500] = 12'b000000_000000;
		Dplus[1501] = 12'b000000_000000;
		Dplus[1502] = 12'b000000_000000;
		Dplus[1503] = 12'b000000_000000;
		Dplus[1504] = 12'b000000_000000;
		Dplus[1505] = 12'b000000_000000;
		Dplus[1506] = 12'b000000_000000;
		Dplus[1507] = 12'b000000_000000;
		Dplus[1508] = 12'b000000_000000;
		Dplus[1509] = 12'b000000_000000;
		Dplus[1510] = 12'b000000_000000;
		Dplus[1511] = 12'b000000_000000;
		Dplus[1512] = 12'b000000_000000;
		Dplus[1513] = 12'b000000_000000;
		Dplus[1514] = 12'b000000_000000;
		Dplus[1515] = 12'b000000_000000;
		Dplus[1516] = 12'b000000_000000;
		Dplus[1517] = 12'b000000_000000;
		Dplus[1518] = 12'b000000_000000;
		Dplus[1519] = 12'b000000_000000;
		Dplus[1520] = 12'b000000_000000;
		Dplus[1521] = 12'b000000_000000;
		Dplus[1522] = 12'b000000_000000;
		Dplus[1523] = 12'b000000_000000;
		Dplus[1524] = 12'b000000_000000;
		Dplus[1525] = 12'b000000_000000;
		Dplus[1526] = 12'b000000_000000;
		Dplus[1527] = 12'b000000_000000;
		Dplus[1528] = 12'b000000_000000;
		Dplus[1529] = 12'b000000_000000;
		Dplus[1530] = 12'b000000_000000;
		Dplus[1531] = 12'b000000_000000;
		Dplus[1532] = 12'b000000_000000;
		Dplus[1533] = 12'b000000_000000;
		Dplus[1534] = 12'b000000_000000;
		Dplus[1535] = 12'b000000_000000;
		Dplus[1536] = 12'b000000_000000;
		Dplus[1537] = 12'b000000_000000;
		Dplus[1538] = 12'b000000_000000;
		Dplus[1539] = 12'b000000_000000;
		Dplus[1540] = 12'b000000_000000;
		Dplus[1541] = 12'b000000_000000;
		Dplus[1542] = 12'b000000_000000;
		Dplus[1543] = 12'b000000_000000;
		Dplus[1544] = 12'b000000_000000;
		Dplus[1545] = 12'b000000_000000;
		Dplus[1546] = 12'b000000_000000;
		Dplus[1547] = 12'b000000_000000;
		Dplus[1548] = 12'b000000_000000;
		Dplus[1549] = 12'b000000_000000;
		Dplus[1550] = 12'b000000_000000;
		Dplus[1551] = 12'b000000_000000;
		Dplus[1552] = 12'b000000_000000;
		Dplus[1553] = 12'b000000_000000;
		Dplus[1554] = 12'b000000_000000;
		Dplus[1555] = 12'b000000_000000;
		Dplus[1556] = 12'b000000_000000;
		Dplus[1557] = 12'b000000_000000;
		Dplus[1558] = 12'b000000_000000;
		Dplus[1559] = 12'b000000_000000;
		Dplus[1560] = 12'b000000_000000;
		Dplus[1561] = 12'b000000_000000;
		Dplus[1562] = 12'b000000_000000;
		Dplus[1563] = 12'b000000_000000;
		Dplus[1564] = 12'b000000_000000;
		Dplus[1565] = 12'b000000_000000;
		Dplus[1566] = 12'b000000_000000;
		Dplus[1567] = 12'b000000_000000;
		Dplus[1568] = 12'b000000_000000;
		Dplus[1569] = 12'b000000_000000;
		Dplus[1570] = 12'b000000_000000;
		Dplus[1571] = 12'b000000_000000;
		Dplus[1572] = 12'b000000_000000;
		Dplus[1573] = 12'b000000_000000;
		Dplus[1574] = 12'b000000_000000;
		Dplus[1575] = 12'b000000_000000;
		Dplus[1576] = 12'b000000_000000;
		Dplus[1577] = 12'b000000_000000;
		Dplus[1578] = 12'b000000_000000;
		Dplus[1579] = 12'b000000_000000;
		Dplus[1580] = 12'b000000_000000;
		Dplus[1581] = 12'b000000_000000;
		Dplus[1582] = 12'b000000_000000;
		Dplus[1583] = 12'b000000_000000;
		Dplus[1584] = 12'b000000_000000;
		Dplus[1585] = 12'b000000_000000;
		Dplus[1586] = 12'b000000_000000;
		Dplus[1587] = 12'b000000_000000;
		Dplus[1588] = 12'b000000_000000;
		Dplus[1589] = 12'b000000_000000;
		Dplus[1590] = 12'b000000_000000;
		Dplus[1591] = 12'b000000_000000;
		Dplus[1592] = 12'b000000_000000;
		Dplus[1593] = 12'b000000_000000;
		Dplus[1594] = 12'b000000_000000;
		Dplus[1595] = 12'b000000_000000;
		Dplus[1596] = 12'b000000_000000;
		Dplus[1597] = 12'b000000_000000;
		Dplus[1598] = 12'b000000_000000;
		Dplus[1599] = 12'b000000_000000;
		Dplus[1600] = 12'b000000_000000;
		Dplus[1601] = 12'b000000_000000;
		Dplus[1602] = 12'b000000_000000;
		Dplus[1603] = 12'b000000_000000;
		Dplus[1604] = 12'b000000_000000;
		Dplus[1605] = 12'b000000_000000;
		Dplus[1606] = 12'b000000_000000;
		Dplus[1607] = 12'b000000_000000;
		Dplus[1608] = 12'b000000_000000;
		Dplus[1609] = 12'b000000_000000;
		Dplus[1610] = 12'b000000_000000;
		Dplus[1611] = 12'b000000_000000;
		Dplus[1612] = 12'b000000_000000;
		Dplus[1613] = 12'b000000_000000;
		Dplus[1614] = 12'b000000_000000;
		Dplus[1615] = 12'b000000_000000;
		Dplus[1616] = 12'b000000_000000;
		Dplus[1617] = 12'b000000_000000;
		Dplus[1618] = 12'b000000_000000;
		Dplus[1619] = 12'b000000_000000;
		Dplus[1620] = 12'b000000_000000;
		Dplus[1621] = 12'b000000_000000;
		Dplus[1622] = 12'b000000_000000;
		Dplus[1623] = 12'b000000_000000;
		Dplus[1624] = 12'b000000_000000;
		Dplus[1625] = 12'b000000_000000;
		Dplus[1626] = 12'b000000_000000;
		Dplus[1627] = 12'b000000_000000;
		Dplus[1628] = 12'b000000_000000;
		Dplus[1629] = 12'b000000_000000;
		Dplus[1630] = 12'b000000_000000;
		Dplus[1631] = 12'b000000_000000;
		Dplus[1632] = 12'b000000_000000;
		Dplus[1633] = 12'b000000_000000;
		Dplus[1634] = 12'b000000_000000;
		Dplus[1635] = 12'b000000_000000;
		Dplus[1636] = 12'b000000_000000;
		Dplus[1637] = 12'b000000_000000;
		Dplus[1638] = 12'b000000_000000;
		Dplus[1639] = 12'b000000_000000;
		Dplus[1640] = 12'b000000_000000;
		Dplus[1641] = 12'b000000_000000;
		Dplus[1642] = 12'b000000_000000;
		Dplus[1643] = 12'b000000_000000;
		Dplus[1644] = 12'b000000_000000;
		Dplus[1645] = 12'b000000_000000;
		Dplus[1646] = 12'b000000_000000;
		Dplus[1647] = 12'b000000_000000;
		Dplus[1648] = 12'b000000_000000;
		Dplus[1649] = 12'b000000_000000;
		Dplus[1650] = 12'b000000_000000;
		Dplus[1651] = 12'b000000_000000;
		Dplus[1652] = 12'b000000_000000;
		Dplus[1653] = 12'b000000_000000;
		Dplus[1654] = 12'b000000_000000;
		Dplus[1655] = 12'b000000_000000;
		Dplus[1656] = 12'b000000_000000;
		Dplus[1657] = 12'b000000_000000;
		Dplus[1658] = 12'b000000_000000;
		Dplus[1659] = 12'b000000_000000;
		Dplus[1660] = 12'b000000_000000;
		Dplus[1661] = 12'b000000_000000;
		Dplus[1662] = 12'b000000_000000;
		Dplus[1663] = 12'b000000_000000;
		Dplus[1664] = 12'b000000_000000;
		Dplus[1665] = 12'b000000_000000;
		Dplus[1666] = 12'b000000_000000;
		Dplus[1667] = 12'b000000_000000;
		Dplus[1668] = 12'b000000_000000;
		Dplus[1669] = 12'b000000_000000;
		Dplus[1670] = 12'b000000_000000;
		Dplus[1671] = 12'b000000_000000;
		Dplus[1672] = 12'b000000_000000;
		Dplus[1673] = 12'b000000_000000;
		Dplus[1674] = 12'b000000_000000;
		Dplus[1675] = 12'b000000_000000;
		Dplus[1676] = 12'b000000_000000;
		Dplus[1677] = 12'b000000_000000;
		Dplus[1678] = 12'b000000_000000;
		Dplus[1679] = 12'b000000_000000;
		Dplus[1680] = 12'b000000_000000;
		Dplus[1681] = 12'b000000_000000;
		Dplus[1682] = 12'b000000_000000;
		Dplus[1683] = 12'b000000_000000;
		Dplus[1684] = 12'b000000_000000;
		Dplus[1685] = 12'b000000_000000;
		Dplus[1686] = 12'b000000_000000;
		Dplus[1687] = 12'b000000_000000;
		Dplus[1688] = 12'b000000_000000;
		Dplus[1689] = 12'b000000_000000;
		Dplus[1690] = 12'b000000_000000;
		Dplus[1691] = 12'b000000_000000;
		Dplus[1692] = 12'b000000_000000;
		Dplus[1693] = 12'b000000_000000;
		Dplus[1694] = 12'b000000_000000;
		Dplus[1695] = 12'b000000_000000;
		Dplus[1696] = 12'b000000_000000;
		Dplus[1697] = 12'b000000_000000;
		Dplus[1698] = 12'b000000_000000;
		Dplus[1699] = 12'b000000_000000;
		Dplus[1700] = 12'b000000_000000;
		Dplus[1701] = 12'b000000_000000;
		Dplus[1702] = 12'b000000_000000;
		Dplus[1703] = 12'b000000_000000;
		Dplus[1704] = 12'b000000_000000;
		Dplus[1705] = 12'b000000_000000;
		Dplus[1706] = 12'b000000_000000;
		Dplus[1707] = 12'b000000_000000;
		Dplus[1708] = 12'b000000_000000;
		Dplus[1709] = 12'b000000_000000;
		Dplus[1710] = 12'b000000_000000;
		Dplus[1711] = 12'b000000_000000;
		Dplus[1712] = 12'b000000_000000;
		Dplus[1713] = 12'b000000_000000;
		Dplus[1714] = 12'b000000_000000;
		Dplus[1715] = 12'b000000_000000;
		Dplus[1716] = 12'b000000_000000;
		Dplus[1717] = 12'b000000_000000;
		Dplus[1718] = 12'b000000_000000;
		Dplus[1719] = 12'b000000_000000;
		Dplus[1720] = 12'b000000_000000;
		Dplus[1721] = 12'b000000_000000;
		Dplus[1722] = 12'b000000_000000;
		Dplus[1723] = 12'b000000_000000;
		Dplus[1724] = 12'b000000_000000;
		Dplus[1725] = 12'b000000_000000;
		Dplus[1726] = 12'b000000_000000;
		Dplus[1727] = 12'b000000_000000;
		Dplus[1728] = 12'b000000_000000;
		Dplus[1729] = 12'b000000_000000;
		Dplus[1730] = 12'b000000_000000;
		Dplus[1731] = 12'b000000_000000;
		Dplus[1732] = 12'b000000_000000;
		Dplus[1733] = 12'b000000_000000;
		Dplus[1734] = 12'b000000_000000;
		Dplus[1735] = 12'b000000_000000;
		Dplus[1736] = 12'b000000_000000;
		Dplus[1737] = 12'b000000_000000;
		Dplus[1738] = 12'b000000_000000;
		Dplus[1739] = 12'b000000_000000;
		Dplus[1740] = 12'b000000_000000;
		Dplus[1741] = 12'b000000_000000;
		Dplus[1742] = 12'b000000_000000;
		Dplus[1743] = 12'b000000_000000;
		Dplus[1744] = 12'b000000_000000;
		Dplus[1745] = 12'b000000_000000;
		Dplus[1746] = 12'b000000_000000;
		Dplus[1747] = 12'b000000_000000;
		Dplus[1748] = 12'b000000_000000;
		Dplus[1749] = 12'b000000_000000;
		Dplus[1750] = 12'b000000_000000;
		Dplus[1751] = 12'b000000_000000;
		Dplus[1752] = 12'b000000_000000;
		Dplus[1753] = 12'b000000_000000;
		Dplus[1754] = 12'b000000_000000;
		Dplus[1755] = 12'b000000_000000;
		Dplus[1756] = 12'b000000_000000;
		Dplus[1757] = 12'b000000_000000;
		Dplus[1758] = 12'b000000_000000;
		Dplus[1759] = 12'b000000_000000;
		Dplus[1760] = 12'b000000_000000;
		Dplus[1761] = 12'b000000_000000;
		Dplus[1762] = 12'b000000_000000;
		Dplus[1763] = 12'b000000_000000;
		Dplus[1764] = 12'b000000_000000;
		Dplus[1765] = 12'b000000_000000;
		Dplus[1766] = 12'b000000_000000;
		Dplus[1767] = 12'b000000_000000;
		Dplus[1768] = 12'b000000_000000;
		Dplus[1769] = 12'b000000_000000;
		Dplus[1770] = 12'b000000_000000;
		Dplus[1771] = 12'b000000_000000;
		Dplus[1772] = 12'b000000_000000;
		Dplus[1773] = 12'b000000_000000;
		Dplus[1774] = 12'b000000_000000;
		Dplus[1775] = 12'b000000_000000;
		Dplus[1776] = 12'b000000_000000;
		Dplus[1777] = 12'b000000_000000;
		Dplus[1778] = 12'b000000_000000;
		Dplus[1779] = 12'b000000_000000;
		Dplus[1780] = 12'b000000_000000;
		Dplus[1781] = 12'b000000_000000;
		Dplus[1782] = 12'b000000_000000;
		Dplus[1783] = 12'b000000_000000;
		Dplus[1784] = 12'b000000_000000;
		Dplus[1785] = 12'b000000_000000;
		Dplus[1786] = 12'b000000_000000;
		Dplus[1787] = 12'b000000_000000;
		Dplus[1788] = 12'b000000_000000;
		Dplus[1789] = 12'b000000_000000;
		Dplus[1790] = 12'b000000_000000;
		Dplus[1791] = 12'b000000_000000;
		Dplus[1792] = 12'b000000_000000;
		Dplus[1793] = 12'b000000_000000;
		Dplus[1794] = 12'b000000_000000;
		Dplus[1795] = 12'b000000_000000;
		Dplus[1796] = 12'b000000_000000;
		Dplus[1797] = 12'b000000_000000;
		Dplus[1798] = 12'b000000_000000;
		Dplus[1799] = 12'b000000_000000;
		Dplus[1800] = 12'b000000_000000;
		Dplus[1801] = 12'b000000_000000;
		Dplus[1802] = 12'b000000_000000;
		Dplus[1803] = 12'b000000_000000;
		Dplus[1804] = 12'b000000_000000;
		Dplus[1805] = 12'b000000_000000;
		Dplus[1806] = 12'b000000_000000;
		Dplus[1807] = 12'b000000_000000;
		Dplus[1808] = 12'b000000_000000;
		Dplus[1809] = 12'b000000_000000;
		Dplus[1810] = 12'b000000_000000;
		Dplus[1811] = 12'b000000_000000;
		Dplus[1812] = 12'b000000_000000;
		Dplus[1813] = 12'b000000_000000;
		Dplus[1814] = 12'b000000_000000;
		Dplus[1815] = 12'b000000_000000;
		Dplus[1816] = 12'b000000_000000;
		Dplus[1817] = 12'b000000_000000;
		Dplus[1818] = 12'b000000_000000;
		Dplus[1819] = 12'b000000_000000;
		Dplus[1820] = 12'b000000_000000;
		Dplus[1821] = 12'b000000_000000;
		Dplus[1822] = 12'b000000_000000;
		Dplus[1823] = 12'b000000_000000;
		Dplus[1824] = 12'b000000_000000;
		Dplus[1825] = 12'b000000_000000;
		Dplus[1826] = 12'b000000_000000;
		Dplus[1827] = 12'b000000_000000;
		Dplus[1828] = 12'b000000_000000;
		Dplus[1829] = 12'b000000_000000;
		Dplus[1830] = 12'b000000_000000;
		Dplus[1831] = 12'b000000_000000;
		Dplus[1832] = 12'b000000_000000;
		Dplus[1833] = 12'b000000_000000;
		Dplus[1834] = 12'b000000_000000;
		Dplus[1835] = 12'b000000_000000;
		Dplus[1836] = 12'b000000_000000;
		Dplus[1837] = 12'b000000_000000;
		Dplus[1838] = 12'b000000_000000;
		Dplus[1839] = 12'b000000_000000;
		Dplus[1840] = 12'b000000_000000;
		Dplus[1841] = 12'b000000_000000;
		Dplus[1842] = 12'b000000_000000;
		Dplus[1843] = 12'b000000_000000;
		Dplus[1844] = 12'b000000_000000;
		Dplus[1845] = 12'b000000_000000;
		Dplus[1846] = 12'b000000_000000;
		Dplus[1847] = 12'b000000_000000;
		Dplus[1848] = 12'b000000_000000;
		Dplus[1849] = 12'b000000_000000;
		Dplus[1850] = 12'b000000_000000;
		Dplus[1851] = 12'b000000_000000;
		Dplus[1852] = 12'b000000_000000;
		Dplus[1853] = 12'b000000_000000;
		Dplus[1854] = 12'b000000_000000;
		Dplus[1855] = 12'b000000_000000;
		Dplus[1856] = 12'b000000_000000;
		Dplus[1857] = 12'b000000_000000;
		Dplus[1858] = 12'b000000_000000;
		Dplus[1859] = 12'b000000_000000;
		Dplus[1860] = 12'b000000_000000;
		Dplus[1861] = 12'b000000_000000;
		Dplus[1862] = 12'b000000_000000;
		Dplus[1863] = 12'b000000_000000;
		Dplus[1864] = 12'b000000_000000;
		Dplus[1865] = 12'b000000_000000;
		Dplus[1866] = 12'b000000_000000;
		Dplus[1867] = 12'b000000_000000;
		Dplus[1868] = 12'b000000_000000;
		Dplus[1869] = 12'b000000_000000;
		Dplus[1870] = 12'b000000_000000;
		Dplus[1871] = 12'b000000_000000;
		Dplus[1872] = 12'b000000_000000;
		Dplus[1873] = 12'b000000_000000;
		Dplus[1874] = 12'b000000_000000;
		Dplus[1875] = 12'b000000_000000;
		Dplus[1876] = 12'b000000_000000;
		Dplus[1877] = 12'b000000_000000;
		Dplus[1878] = 12'b000000_000000;
		Dplus[1879] = 12'b000000_000000;
		Dplus[1880] = 12'b000000_000000;
		Dplus[1881] = 12'b000000_000000;
		Dplus[1882] = 12'b000000_000000;
		Dplus[1883] = 12'b000000_000000;
		Dplus[1884] = 12'b000000_000000;
		Dplus[1885] = 12'b000000_000000;
		Dplus[1886] = 12'b000000_000000;
		Dplus[1887] = 12'b000000_000000;
		Dplus[1888] = 12'b000000_000000;
		Dplus[1889] = 12'b000000_000000;
		Dplus[1890] = 12'b000000_000000;
		Dplus[1891] = 12'b000000_000000;
		Dplus[1892] = 12'b000000_000000;
		Dplus[1893] = 12'b000000_000000;
		Dplus[1894] = 12'b000000_000000;
		Dplus[1895] = 12'b000000_000000;
		Dplus[1896] = 12'b000000_000000;
		Dplus[1897] = 12'b000000_000000;
		Dplus[1898] = 12'b000000_000000;
		Dplus[1899] = 12'b000000_000000;
		Dplus[1900] = 12'b000000_000000;
		Dplus[1901] = 12'b000000_000000;
		Dplus[1902] = 12'b000000_000000;
		Dplus[1903] = 12'b000000_000000;
		Dplus[1904] = 12'b000000_000000;
		Dplus[1905] = 12'b000000_000000;
		Dplus[1906] = 12'b000000_000000;
		Dplus[1907] = 12'b000000_000000;
		Dplus[1908] = 12'b000000_000000;
		Dplus[1909] = 12'b000000_000000;
		Dplus[1910] = 12'b000000_000000;
		Dplus[1911] = 12'b000000_000000;
		Dplus[1912] = 12'b000000_000000;
		Dplus[1913] = 12'b000000_000000;
		Dplus[1914] = 12'b000000_000000;
		Dplus[1915] = 12'b000000_000000;
		Dplus[1916] = 12'b000000_000000;
		Dplus[1917] = 12'b000000_000000;
		Dplus[1918] = 12'b000000_000000;
		Dplus[1919] = 12'b000000_000000;
		Dplus[1920] = 12'b000000_000000;
		Dplus[1921] = 12'b000000_000000;
		Dplus[1922] = 12'b000000_000000;
		Dplus[1923] = 12'b000000_000000;
		Dplus[1924] = 12'b000000_000000;
		Dplus[1925] = 12'b000000_000000;
		Dplus[1926] = 12'b000000_000000;
		Dplus[1927] = 12'b000000_000000;
		Dplus[1928] = 12'b000000_000000;
		Dplus[1929] = 12'b000000_000000;
		Dplus[1930] = 12'b000000_000000;
		Dplus[1931] = 12'b000000_000000;
		Dplus[1932] = 12'b000000_000000;
		Dplus[1933] = 12'b000000_000000;
		Dplus[1934] = 12'b000000_000000;
		Dplus[1935] = 12'b000000_000000;
		Dplus[1936] = 12'b000000_000000;
		Dplus[1937] = 12'b000000_000000;
		Dplus[1938] = 12'b000000_000000;
		Dplus[1939] = 12'b000000_000000;
		Dplus[1940] = 12'b000000_000000;
		Dplus[1941] = 12'b000000_000000;
		Dplus[1942] = 12'b000000_000000;
		Dplus[1943] = 12'b000000_000000;
		Dplus[1944] = 12'b000000_000000;
		Dplus[1945] = 12'b000000_000000;
		Dplus[1946] = 12'b000000_000000;
		Dplus[1947] = 12'b000000_000000;
		Dplus[1948] = 12'b000000_000000;
		Dplus[1949] = 12'b000000_000000;
		Dplus[1950] = 12'b000000_000000;
		Dplus[1951] = 12'b000000_000000;
		Dplus[1952] = 12'b000000_000000;
		Dplus[1953] = 12'b000000_000000;
		Dplus[1954] = 12'b000000_000000;
		Dplus[1955] = 12'b000000_000000;
		Dplus[1956] = 12'b000000_000000;
		Dplus[1957] = 12'b000000_000000;
		Dplus[1958] = 12'b000000_000000;
		Dplus[1959] = 12'b000000_000000;
		Dplus[1960] = 12'b000000_000000;
		Dplus[1961] = 12'b000000_000000;
		Dplus[1962] = 12'b000000_000000;
		Dplus[1963] = 12'b000000_000000;
		Dplus[1964] = 12'b000000_000000;
		Dplus[1965] = 12'b000000_000000;
		Dplus[1966] = 12'b000000_000000;
		Dplus[1967] = 12'b000000_000000;
		Dplus[1968] = 12'b000000_000000;
		Dplus[1969] = 12'b000000_000000;
		Dplus[1970] = 12'b000000_000000;
		Dplus[1971] = 12'b000000_000000;
		Dplus[1972] = 12'b000000_000000;
		Dplus[1973] = 12'b000000_000000;
		Dplus[1974] = 12'b000000_000000;
		Dplus[1975] = 12'b000000_000000;
		Dplus[1976] = 12'b000000_000000;
		Dplus[1977] = 12'b000000_000000;
		Dplus[1978] = 12'b000000_000000;
		Dplus[1979] = 12'b000000_000000;
		Dplus[1980] = 12'b000000_000000;
		Dplus[1981] = 12'b000000_000000;
		Dplus[1982] = 12'b000000_000000;
		Dplus[1983] = 12'b000000_000000;
		Dplus[1984] = 12'b000000_000000;
		Dplus[1985] = 12'b000000_000000;
		Dplus[1986] = 12'b000000_000000;
		Dplus[1987] = 12'b000000_000000;
		Dplus[1988] = 12'b000000_000000;
		Dplus[1989] = 12'b000000_000000;
		Dplus[1990] = 12'b000000_000000;
		Dplus[1991] = 12'b000000_000000;
		Dplus[1992] = 12'b000000_000000;
		Dplus[1993] = 12'b000000_000000;
		Dplus[1994] = 12'b000000_000000;
		Dplus[1995] = 12'b000000_000000;
		Dplus[1996] = 12'b000000_000000;
		Dplus[1997] = 12'b000000_000000;
		Dplus[1998] = 12'b000000_000000;
		Dplus[1999] = 12'b000000_000000;
		Dplus[2000] = 12'b000000_000000;
		Dplus[2001] = 12'b000000_000000;
		Dplus[2002] = 12'b000000_000000;
		Dplus[2003] = 12'b000000_000000;
		Dplus[2004] = 12'b000000_000000;
		Dplus[2005] = 12'b000000_000000;
		Dplus[2006] = 12'b000000_000000;
		Dplus[2007] = 12'b000000_000000;
		Dplus[2008] = 12'b000000_000000;
		Dplus[2009] = 12'b000000_000000;
		Dplus[2010] = 12'b000000_000000;
		Dplus[2011] = 12'b000000_000000;
		Dplus[2012] = 12'b000000_000000;
		Dplus[2013] = 12'b000000_000000;
		Dplus[2014] = 12'b000000_000000;
		Dplus[2015] = 12'b000000_000000;
		Dplus[2016] = 12'b000000_000000;
		Dplus[2017] = 12'b000000_000000;
		Dplus[2018] = 12'b000000_000000;
		Dplus[2019] = 12'b000000_000000;
		Dplus[2020] = 12'b000000_000000;
		Dplus[2021] = 12'b000000_000000;
		Dplus[2022] = 12'b000000_000000;
		Dplus[2023] = 12'b000000_000000;
		Dplus[2024] = 12'b000000_000000;
		Dplus[2025] = 12'b000000_000000;
		Dplus[2026] = 12'b000000_000000;
		Dplus[2027] = 12'b000000_000000;
		Dplus[2028] = 12'b000000_000000;
		Dplus[2029] = 12'b000000_000000;
		Dplus[2030] = 12'b000000_000000;
		Dplus[2031] = 12'b000000_000000;
		Dplus[2032] = 12'b000000_000000;
		Dplus[2033] = 12'b000000_000000;
		Dplus[2034] = 12'b000000_000000;
		Dplus[2035] = 12'b000000_000000;
		Dplus[2036] = 12'b000000_000000;
		Dplus[2037] = 12'b000000_000000;
		Dplus[2038] = 12'b000000_000000;
		Dplus[2039] = 12'b000000_000000;
		Dplus[2040] = 12'b000000_000000;
		Dplus[2041] = 12'b000000_000000;
		Dplus[2042] = 12'b000000_000000;
		Dplus[2043] = 12'b000000_000000;
		Dplus[2044] = 12'b000000_000000;
		Dplus[2045] = 12'b000000_000000;
		Dplus[2046] = 12'b000000_000000;
		Dplus[2047] = 12'b000000_000000;
end
endmodule
