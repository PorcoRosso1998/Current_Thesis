module Tables();
	reg [11:0] Dplus[127:0];
	reg [11:0] Dminus[127:0];
	reg [5:0] DminusInteger[31:0];
	reg [5:0] DplusInteger[31:0];
	initial begin
		Dminus[1] = 12'b111001_011110;
		Dminus[2] = 12'b111010_011101;
		Dminus[3] = 12'b111011_000010;
		Dminus[4] = 12'b111011_011100;
		Dminus[5] = 12'b111011_110000;
		Dminus[6] = 12'b111100_000001;
		Dminus[7] = 12'b111100_001110;
		Dminus[8] = 12'b111100_011010;
		Dminus[9] = 12'b111100_100101;
		Dminus[10] = 12'b111100_101110;
		Dminus[11] = 12'b111100_110110;
		Dminus[12] = 12'b111100_111110;
		Dminus[13] = 12'b111101_000101;
		Dminus[14] = 12'b111101_001011;
		Dminus[15] = 12'b111101_010001;
		Dminus[16] = 12'b111101_010110;
		Dminus[17] = 12'b111101_011011;
		Dminus[18] = 12'b111101_100000;
		Dminus[19] = 12'b111101_100101;
		Dminus[20] = 12'b111101_101001;
		Dminus[21] = 12'b111101_101101;
		Dminus[22] = 12'b111101_110001;
		Dminus[23] = 12'b111101_110100;
		Dminus[24] = 12'b111101_111000;
		Dminus[25] = 12'b111101_111011;
		Dminus[26] = 12'b111101_111110;
		Dminus[27] = 12'b111110_000001;
		Dminus[28] = 12'b111110_000100;
		Dminus[29] = 12'b111110_000111;
		Dminus[30] = 12'b111110_001010;
		Dminus[31] = 12'b111110_001100;
		Dminus[32] = 12'b111110_001111;
		Dminus[33] = 12'b111110_010001;
		Dminus[34] = 12'b111110_010011;
		Dminus[35] = 12'b111110_010101;
		Dminus[36] = 12'b111110_011000;
		Dminus[37] = 12'b111110_011010;
		Dminus[38] = 12'b111110_011100;
		Dminus[39] = 12'b111110_011110;
		Dminus[40] = 12'b111110_011111;
		Dminus[41] = 12'b111110_100001;
		Dminus[42] = 12'b111110_100011;
		Dminus[43] = 12'b111110_100101;
		Dminus[44] = 12'b111110_100110;
		Dminus[45] = 12'b111110_101000;
		Dminus[46] = 12'b111110_101010;
		Dminus[47] = 12'b111110_101011;
		Dminus[48] = 12'b111110_101101;
		Dminus[49] = 12'b111110_101110;
		Dminus[50] = 12'b111110_101111;
		Dminus[51] = 12'b111110_110001;
		Dminus[52] = 12'b111110_110010;
		Dminus[53] = 12'b111110_110100;
		Dminus[54] = 12'b111110_110101;
		Dminus[55] = 12'b111110_110110;
		Dminus[56] = 12'b111110_110111;
		Dminus[57] = 12'b111110_111000;
		Dminus[58] = 12'b111110_111010;
		Dminus[59] = 12'b111110_111011;
		Dminus[60] = 12'b111110_111100;
		Dminus[61] = 12'b111110_111101;
		Dminus[62] = 12'b111110_111110;
		Dminus[63] = 12'b111110_111111;
		Dminus[64] = 12'b111111_000000;
		Dminus[65] = 12'b111111_000001;
		Dminus[66] = 12'b111111_000010;
		Dminus[67] = 12'b111111_000011;
		Dminus[68] = 12'b111111_000100;
		Dminus[69] = 12'b111111_000101;
		Dminus[70] = 12'b111111_000110;
		Dminus[71] = 12'b111111_000111;
		Dminus[72] = 12'b111111_000111;
		Dminus[73] = 12'b111111_001000;
		Dminus[74] = 12'b111111_001001;
		Dminus[75] = 12'b111111_001010;
		Dminus[76] = 12'b111111_001011;
		Dminus[77] = 12'b111111_001011;
		Dminus[78] = 12'b111111_001100;
		Dminus[79] = 12'b111111_001101;
		Dminus[80] = 12'b111111_001110;
		Dminus[81] = 12'b111111_001110;
		Dminus[82] = 12'b111111_001111;
		Dminus[83] = 12'b111111_010000;
		Dminus[84] = 12'b111111_010000;
		Dminus[85] = 12'b111111_010001;
		Dminus[86] = 12'b111111_010010;
		Dminus[87] = 12'b111111_010010;
		Dminus[88] = 12'b111111_010011;
		Dminus[89] = 12'b111111_010100;
		Dminus[90] = 12'b111111_010100;
		Dminus[91] = 12'b111111_010101;
		Dminus[92] = 12'b111111_010101;
		Dminus[93] = 12'b111111_010110;
		Dminus[94] = 12'b111111_010111;
		Dminus[95] = 12'b111111_010111;
		Dminus[96] = 12'b111111_011000;
		Dminus[97] = 12'b111111_011000;
		Dminus[98] = 12'b111111_011001;
		Dminus[99] = 12'b111111_011001;
		Dminus[100] = 12'b111111_011010;
		Dminus[101] = 12'b111111_011010;
		Dminus[102] = 12'b111111_011011;
		Dminus[103] = 12'b111111_011011;
		Dminus[104] = 12'b111111_011100;
		Dminus[105] = 12'b111111_011100;
		Dminus[106] = 12'b111111_011101;
		Dminus[107] = 12'b111111_011101;
		Dminus[108] = 12'b111111_011110;
		Dminus[109] = 12'b111111_011110;
		Dminus[110] = 12'b111111_011111;
		Dminus[111] = 12'b111111_011111;
		Dminus[112] = 12'b111111_011111;
		Dminus[113] = 12'b111111_100000;
		Dminus[114] = 12'b111111_100000;
		Dminus[115] = 12'b111111_100001;
		Dminus[116] = 12'b111111_100001;
		Dminus[117] = 12'b111111_100001;
		Dminus[118] = 12'b111111_100010;
		Dminus[119] = 12'b111111_100010;
		Dminus[120] = 12'b111111_100011;
		Dminus[121] = 12'b111111_100011;
		Dminus[122] = 12'b111111_100011;
		Dminus[123] = 12'b111111_100100;
		Dminus[124] = 12'b111111_100100;
		Dminus[125] = 12'b111111_100100;
		Dminus[126] = 12'b111111_100101;
		Dminus[127] = 12'b111111_100101;
		Dplus[1] = 12'b000001_000000;
		Dplus[2] = 12'b000000_111111;
		Dplus[3] = 12'b000000_111111;
		Dplus[4] = 12'b000000_111110;
		Dplus[5] = 12'b000000_111110;
		Dplus[6] = 12'b000000_111101;
		Dplus[7] = 12'b000000_111101;
		Dplus[8] = 12'b000000_111100;
		Dplus[9] = 12'b000000_111100;
		Dplus[10] = 12'b000000_111011;
		Dplus[11] = 12'b000000_111011;
		Dplus[12] = 12'b000000_111010;
		Dplus[13] = 12'b000000_111010;
		Dplus[14] = 12'b000000_111001;
		Dplus[15] = 12'b000000_111001;
		Dplus[16] = 12'b000000_111000;
		Dplus[17] = 12'b000000_111000;
		Dplus[18] = 12'b000000_110111;
		Dplus[19] = 12'b000000_110111;
		Dplus[20] = 12'b000000_110111;
		Dplus[21] = 12'b000000_110110;
		Dplus[22] = 12'b000000_110110;
		Dplus[23] = 12'b000000_110101;
		Dplus[24] = 12'b000000_110101;
		Dplus[25] = 12'b000000_110100;
		Dplus[26] = 12'b000000_110100;
		Dplus[27] = 12'b000000_110011;
		Dplus[28] = 12'b000000_110011;
		Dplus[29] = 12'b000000_110011;
		Dplus[30] = 12'b000000_110010;
		Dplus[31] = 12'b000000_110010;
		Dplus[32] = 12'b000000_110001;
		Dplus[33] = 12'b000000_110001;
		Dplus[34] = 12'b000000_110001;
		Dplus[35] = 12'b000000_110000;
		Dplus[36] = 12'b000000_110000;
		Dplus[37] = 12'b000000_101111;
		Dplus[38] = 12'b000000_101111;
		Dplus[39] = 12'b000000_101111;
		Dplus[40] = 12'b000000_101110;
		Dplus[41] = 12'b000000_101110;
		Dplus[42] = 12'b000000_101101;
		Dplus[43] = 12'b000000_101101;
		Dplus[44] = 12'b000000_101101;
		Dplus[45] = 12'b000000_101100;
		Dplus[46] = 12'b000000_101100;
		Dplus[47] = 12'b000000_101011;
		Dplus[48] = 12'b000000_101011;
		Dplus[49] = 12'b000000_101011;
		Dplus[50] = 12'b000000_101010;
		Dplus[51] = 12'b000000_101010;
		Dplus[52] = 12'b000000_101010;
		Dplus[53] = 12'b000000_101001;
		Dplus[54] = 12'b000000_101001;
		Dplus[55] = 12'b000000_101001;
		Dplus[56] = 12'b000000_101000;
		Dplus[57] = 12'b000000_101000;
		Dplus[58] = 12'b000000_100111;
		Dplus[59] = 12'b000000_100111;
		Dplus[60] = 12'b000000_100111;
		Dplus[61] = 12'b000000_100110;
		Dplus[62] = 12'b000000_100110;
		Dplus[63] = 12'b000000_100110;
		Dplus[64] = 12'b000000_100101;
		Dplus[65] = 12'b000000_100101;
		Dplus[66] = 12'b000000_100101;
		Dplus[67] = 12'b000000_100100;
		Dplus[68] = 12'b000000_100100;
		Dplus[69] = 12'b000000_100100;
		Dplus[70] = 12'b000000_100011;
		Dplus[71] = 12'b000000_100011;
		Dplus[72] = 12'b000000_100011;
		Dplus[73] = 12'b000000_100011;
		Dplus[74] = 12'b000000_100010;
		Dplus[75] = 12'b000000_100010;
		Dplus[76] = 12'b000000_100010;
		Dplus[77] = 12'b000000_100001;
		Dplus[78] = 12'b000000_100001;
		Dplus[79] = 12'b000000_100001;
		Dplus[80] = 12'b000000_100000;
		Dplus[81] = 12'b000000_100000;
		Dplus[82] = 12'b000000_100000;
		Dplus[83] = 12'b000000_100000;
		Dplus[84] = 12'b000000_011111;
		Dplus[85] = 12'b000000_011111;
		Dplus[86] = 12'b000000_011111;
		Dplus[87] = 12'b000000_011110;
		Dplus[88] = 12'b000000_011110;
		Dplus[89] = 12'b000000_011110;
		Dplus[90] = 12'b000000_011110;
		Dplus[91] = 12'b000000_011101;
		Dplus[92] = 12'b000000_011101;
		Dplus[93] = 12'b000000_011101;
		Dplus[94] = 12'b000000_011100;
		Dplus[95] = 12'b000000_011100;
		Dplus[96] = 12'b000000_011100;
		Dplus[97] = 12'b000000_011100;
		Dplus[98] = 12'b000000_011011;
		Dplus[99] = 12'b000000_011011;
		Dplus[100] = 12'b000000_011011;
		Dplus[101] = 12'b000000_011011;
		Dplus[102] = 12'b000000_011010;
		Dplus[103] = 12'b000000_011010;
		Dplus[104] = 12'b000000_011010;
		Dplus[105] = 12'b000000_011010;
		Dplus[106] = 12'b000000_011001;
		Dplus[107] = 12'b000000_011001;
		Dplus[108] = 12'b000000_011001;
		Dplus[109] = 12'b000000_011001;
		Dplus[110] = 12'b000000_011000;
		Dplus[111] = 12'b000000_011000;
		Dplus[112] = 12'b000000_011000;
		Dplus[113] = 12'b000000_011000;
		Dplus[114] = 12'b000000_011000;
		Dplus[115] = 12'b000000_010111;
		Dplus[116] = 12'b000000_010111;
		Dplus[117] = 12'b000000_010111;
		Dplus[118] = 12'b000000_010111;
		Dplus[119] = 12'b000000_010110;
		Dplus[120] = 12'b000000_010110;
		Dplus[121] = 12'b000000_010110;
		Dplus[122] = 12'b000000_010110;
		Dplus[123] = 12'b000000_010110;
		Dplus[124] = 12'b000000_010101;
		Dplus[125] = 12'b000000_010101;
		Dplus[126] = 12'b000000_010101;
		Dplus[127] = 12'b000000_010101;
		DplusInteger[2] = 12'b000000_010101;
		DplusInteger[3] = 12'b000000_001011;
		DplusInteger[4] = 12'b000000_000110;
		DplusInteger[5] = 12'b000000_000011;
		DplusInteger[6] = 12'b000000_000001;
		DplusInteger[7] = 12'b000000_000001;
		DplusInteger[8] = 12'b000000_000000;
		DplusInteger[9] = 12'b000000_000000;
		DplusInteger[10] = 12'b000000_000000;
		DplusInteger[11] = 12'b000000_000000;
		DplusInteger[12] = 12'b000000_000000;
		DplusInteger[13] = 12'b000000_000000;
		DplusInteger[14] = 12'b000000_000000;
		DplusInteger[15] = 12'b000000_000000;
		DplusInteger[16] = 12'b000000_000000;
		DplusInteger[17] = 12'b000000_000000;
		DplusInteger[18] = 12'b000000_000000;
		DplusInteger[19] = 12'b000000_000000;
		DplusInteger[20] = 12'b000000_000000;
		DplusInteger[21] = 12'b000000_000000;
		DplusInteger[22] = 12'b000000_000000;
		DplusInteger[23] = 12'b000000_000000;
		DplusInteger[24] = 12'b000000_000000;
		DplusInteger[25] = 12'b000000_000000;
		DplusInteger[26] = 12'b000000_000000;
		DplusInteger[27] = 12'b000000_000000;
		DplusInteger[28] = 12'b000000_000000;
		DplusInteger[29] = 12'b000000_000000;
		DplusInteger[30] = 12'b000000_000000;
		DplusInteger[31] = 12'b000000_000000;
		DminusInteger[2] = 12'b111111_100101;
		DminusInteger[3] = 12'b111111_110100;
		DminusInteger[4] = 12'b111111_111010;
		DminusInteger[5] = 12'b111111_111101;
		DminusInteger[6] = 12'b111111_111111;
		DminusInteger[7] = 12'b111111_111111;
		DminusInteger[8] = 12'b000000_000000;
		DminusInteger[9] = 12'b000000_000000;
		DminusInteger[10] = 12'b000000_000000;
		DminusInteger[11] = 12'b000000_000000;
		DminusInteger[12] = 12'b000000_000000;
		DminusInteger[13] = 12'b000000_000000;
		DminusInteger[14] = 12'b000000_000000;
		DminusInteger[15] = 12'b000000_000000;
		DminusInteger[16] = 12'b000000_000000;
		DminusInteger[17] = 12'b000000_000000;
		DminusInteger[18] = 12'b000000_000000;
		DminusInteger[19] = 12'b000000_000000;
		DminusInteger[20] = 12'b000000_000000;
		DminusInteger[21] = 12'b000000_000000;
		DminusInteger[22] = 12'b000000_000000;
		DminusInteger[23] = 12'b000000_000000;
		DminusInteger[24] = 12'b000000_000000;
		DminusInteger[25] = 12'b000000_000000;
		DminusInteger[26] = 12'b000000_000000;
		DminusInteger[27] = 12'b000000_000000;
		DminusInteger[28] = 12'b000000_000000;
		DminusInteger[29] = 12'b000000_000000;
		DminusInteger[30] = 12'b000000_000000;
		DminusInteger[31] = 12'b000000_000000;
end
endmodule
