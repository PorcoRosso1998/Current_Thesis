module Tables();
	reg [17:0] Dplus[1023:0];
	reg [17:0] Dminus[1023:0];
	reg [17:0] DminusInteger[255:0];
	reg [17:0] DplusInteger[255:0];
	initial begin
		Dminus[1] = 18'b111110110_011110001;
		Dminus[2] = 18'b111110111_011110000;
		Dminus[3] = 18'b111111000_000011011;
		Dminus[4] = 18'b111111000_011101111;
		Dminus[5] = 18'b111111000_110010100;
		Dminus[6] = 18'b111111001_000011010;
		Dminus[7] = 18'b111111001_010001011;
		Dminus[8] = 18'b111111001_011101101;
		Dminus[9] = 18'b111111001_101000100;
		Dminus[10] = 18'b111111001_110010001;
		Dminus[11] = 18'b111111001_111010111;
		Dminus[12] = 18'b111111010_000010111;
		Dminus[13] = 18'b111111010_001010001;
		Dminus[14] = 18'b111111010_010001000;
		Dminus[15] = 18'b111111010_010111010;
		Dminus[16] = 18'b111111010_011101001;
		Dminus[17] = 18'b111111010_100010110;
		Dminus[18] = 18'b111111010_100111111;
		Dminus[19] = 18'b111111010_101100111;
		Dminus[20] = 18'b111111010_110001100;
		Dminus[21] = 18'b111111010_110110000;
		Dminus[22] = 18'b111111010_111010010;
		Dminus[23] = 18'b111111010_111110010;
		Dminus[24] = 18'b111111011_000010001;
		Dminus[25] = 18'b111111011_000101110;
		Dminus[26] = 18'b111111011_001001011;
		Dminus[27] = 18'b111111011_001100110;
		Dminus[28] = 18'b111111011_010000001;
		Dminus[29] = 18'b111111011_010011010;
		Dminus[30] = 18'b111111011_010110011;
		Dminus[31] = 18'b111111011_011001010;
		Dminus[32] = 18'b111111011_011100001;
		Dminus[33] = 18'b111111011_011111000;
		Dminus[34] = 18'b111111011_100001101;
		Dminus[35] = 18'b111111011_100100010;
		Dminus[36] = 18'b111111011_100110110;
		Dminus[37] = 18'b111111011_101001010;
		Dminus[38] = 18'b111111011_101011101;
		Dminus[39] = 18'b111111011_101110000;
		Dminus[40] = 18'b111111011_110000010;
		Dminus[41] = 18'b111111011_110010100;
		Dminus[42] = 18'b111111011_110100101;
		Dminus[43] = 18'b111111011_110110110;
		Dminus[44] = 18'b111111011_111000111;
		Dminus[45] = 18'b111111011_111010111;
		Dminus[46] = 18'b111111011_111100110;
		Dminus[47] = 18'b111111011_111110110;
		Dminus[48] = 18'b111111100_000000101;
		Dminus[49] = 18'b111111100_000010100;
		Dminus[50] = 18'b111111100_000100010;
		Dminus[51] = 18'b111111100_000110000;
		Dminus[52] = 18'b111111100_000111110;
		Dminus[53] = 18'b111111100_001001100;
		Dminus[54] = 18'b111111100_001011001;
		Dminus[55] = 18'b111111100_001100110;
		Dminus[56] = 18'b111111100_001110011;
		Dminus[57] = 18'b111111100_001111111;
		Dminus[58] = 18'b111111100_010001100;
		Dminus[59] = 18'b111111100_010011000;
		Dminus[60] = 18'b111111100_010100100;
		Dminus[61] = 18'b111111100_010110000;
		Dminus[62] = 18'b111111100_010111011;
		Dminus[63] = 18'b111111100_011000110;
		Dminus[64] = 18'b111111100_011010010;
		Dminus[65] = 18'b111111100_011011100;
		Dminus[66] = 18'b111111100_011100111;
		Dminus[67] = 18'b111111100_011110010;
		Dminus[68] = 18'b111111100_011111100;
		Dminus[69] = 18'b111111100_100000111;
		Dminus[70] = 18'b111111100_100010001;
		Dminus[71] = 18'b111111100_100011011;
		Dminus[72] = 18'b111111100_100100101;
		Dminus[73] = 18'b111111100_100101110;
		Dminus[74] = 18'b111111100_100111000;
		Dminus[75] = 18'b111111100_101000001;
		Dminus[76] = 18'b111111100_101001011;
		Dminus[77] = 18'b111111100_101010100;
		Dminus[78] = 18'b111111100_101011101;
		Dminus[79] = 18'b111111100_101100110;
		Dminus[80] = 18'b111111100_101101110;
		Dminus[81] = 18'b111111100_101110111;
		Dminus[82] = 18'b111111100_110000000;
		Dminus[83] = 18'b111111100_110001000;
		Dminus[84] = 18'b111111100_110010001;
		Dminus[85] = 18'b111111100_110011001;
		Dminus[86] = 18'b111111100_110100001;
		Dminus[87] = 18'b111111100_110101001;
		Dminus[88] = 18'b111111100_110110001;
		Dminus[89] = 18'b111111100_110111001;
		Dminus[90] = 18'b111111100_111000001;
		Dminus[91] = 18'b111111100_111001000;
		Dminus[92] = 18'b111111100_111010000;
		Dminus[93] = 18'b111111100_111010111;
		Dminus[94] = 18'b111111100_111011111;
		Dminus[95] = 18'b111111100_111100110;
		Dminus[96] = 18'b111111100_111101101;
		Dminus[97] = 18'b111111100_111110100;
		Dminus[98] = 18'b111111100_111111100;
		Dminus[99] = 18'b111111101_000000011;
		Dminus[100] = 18'b111111101_000001001;
		Dminus[101] = 18'b111111101_000010000;
		Dminus[102] = 18'b111111101_000010111;
		Dminus[103] = 18'b111111101_000011110;
		Dminus[104] = 18'b111111101_000100101;
		Dminus[105] = 18'b111111101_000101011;
		Dminus[106] = 18'b111111101_000110010;
		Dminus[107] = 18'b111111101_000111000;
		Dminus[108] = 18'b111111101_000111110;
		Dminus[109] = 18'b111111101_001000101;
		Dminus[110] = 18'b111111101_001001011;
		Dminus[111] = 18'b111111101_001010001;
		Dminus[112] = 18'b111111101_001010111;
		Dminus[113] = 18'b111111101_001011101;
		Dminus[114] = 18'b111111101_001100011;
		Dminus[115] = 18'b111111101_001101001;
		Dminus[116] = 18'b111111101_001101111;
		Dminus[117] = 18'b111111101_001110101;
		Dminus[118] = 18'b111111101_001111011;
		Dminus[119] = 18'b111111101_010000001;
		Dminus[120] = 18'b111111101_010000110;
		Dminus[121] = 18'b111111101_010001100;
		Dminus[122] = 18'b111111101_010010010;
		Dminus[123] = 18'b111111101_010010111;
		Dminus[124] = 18'b111111101_010011101;
		Dminus[125] = 18'b111111101_010100010;
		Dminus[126] = 18'b111111101_010101000;
		Dminus[127] = 18'b111111101_010101101;
		Dminus[128] = 18'b111111101_010110010;
		Dminus[129] = 18'b111111101_010110111;
		Dminus[130] = 18'b111111101_010111101;
		Dminus[131] = 18'b111111101_011000010;
		Dminus[132] = 18'b111111101_011000111;
		Dminus[133] = 18'b111111101_011001100;
		Dminus[134] = 18'b111111101_011010001;
		Dminus[135] = 18'b111111101_011010110;
		Dminus[136] = 18'b111111101_011011011;
		Dminus[137] = 18'b111111101_011100000;
		Dminus[138] = 18'b111111101_011100101;
		Dminus[139] = 18'b111111101_011101010;
		Dminus[140] = 18'b111111101_011101111;
		Dminus[141] = 18'b111111101_011110011;
		Dminus[142] = 18'b111111101_011111000;
		Dminus[143] = 18'b111111101_011111101;
		Dminus[144] = 18'b111111101_100000001;
		Dminus[145] = 18'b111111101_100000110;
		Dminus[146] = 18'b111111101_100001011;
		Dminus[147] = 18'b111111101_100001111;
		Dminus[148] = 18'b111111101_100010100;
		Dminus[149] = 18'b111111101_100011000;
		Dminus[150] = 18'b111111101_100011101;
		Dminus[151] = 18'b111111101_100100001;
		Dminus[152] = 18'b111111101_100100110;
		Dminus[153] = 18'b111111101_100101010;
		Dminus[154] = 18'b111111101_100101110;
		Dminus[155] = 18'b111111101_100110011;
		Dminus[156] = 18'b111111101_100110111;
		Dminus[157] = 18'b111111101_100111011;
		Dminus[158] = 18'b111111101_100111111;
		Dminus[159] = 18'b111111101_101000011;
		Dminus[160] = 18'b111111101_101001000;
		Dminus[161] = 18'b111111101_101001100;
		Dminus[162] = 18'b111111101_101010000;
		Dminus[163] = 18'b111111101_101010100;
		Dminus[164] = 18'b111111101_101011000;
		Dminus[165] = 18'b111111101_101011100;
		Dminus[166] = 18'b111111101_101100000;
		Dminus[167] = 18'b111111101_101100100;
		Dminus[168] = 18'b111111101_101101000;
		Dminus[169] = 18'b111111101_101101100;
		Dminus[170] = 18'b111111101_101110000;
		Dminus[171] = 18'b111111101_101110011;
		Dminus[172] = 18'b111111101_101110111;
		Dminus[173] = 18'b111111101_101111011;
		Dminus[174] = 18'b111111101_101111111;
		Dminus[175] = 18'b111111101_110000011;
		Dminus[176] = 18'b111111101_110000110;
		Dminus[177] = 18'b111111101_110001010;
		Dminus[178] = 18'b111111101_110001110;
		Dminus[179] = 18'b111111101_110010001;
		Dminus[180] = 18'b111111101_110010101;
		Dminus[181] = 18'b111111101_110011001;
		Dminus[182] = 18'b111111101_110011100;
		Dminus[183] = 18'b111111101_110100000;
		Dminus[184] = 18'b111111101_110100011;
		Dminus[185] = 18'b111111101_110100111;
		Dminus[186] = 18'b111111101_110101010;
		Dminus[187] = 18'b111111101_110101110;
		Dminus[188] = 18'b111111101_110110001;
		Dminus[189] = 18'b111111101_110110101;
		Dminus[190] = 18'b111111101_110111000;
		Dminus[191] = 18'b111111101_110111011;
		Dminus[192] = 18'b111111101_110111111;
		Dminus[193] = 18'b111111101_111000010;
		Dminus[194] = 18'b111111101_111000110;
		Dminus[195] = 18'b111111101_111001001;
		Dminus[196] = 18'b111111101_111001100;
		Dminus[197] = 18'b111111101_111001111;
		Dminus[198] = 18'b111111101_111010011;
		Dminus[199] = 18'b111111101_111010110;
		Dminus[200] = 18'b111111101_111011001;
		Dminus[201] = 18'b111111101_111011100;
		Dminus[202] = 18'b111111101_111100000;
		Dminus[203] = 18'b111111101_111100011;
		Dminus[204] = 18'b111111101_111100110;
		Dminus[205] = 18'b111111101_111101001;
		Dminus[206] = 18'b111111101_111101100;
		Dminus[207] = 18'b111111101_111101111;
		Dminus[208] = 18'b111111101_111110010;
		Dminus[209] = 18'b111111101_111110101;
		Dminus[210] = 18'b111111101_111111000;
		Dminus[211] = 18'b111111101_111111011;
		Dminus[212] = 18'b111111101_111111111;
		Dminus[213] = 18'b111111110_000000010;
		Dminus[214] = 18'b111111110_000000100;
		Dminus[215] = 18'b111111110_000000111;
		Dminus[216] = 18'b111111110_000001010;
		Dminus[217] = 18'b111111110_000001101;
		Dminus[218] = 18'b111111110_000010000;
		Dminus[219] = 18'b111111110_000010011;
		Dminus[220] = 18'b111111110_000010110;
		Dminus[221] = 18'b111111110_000011001;
		Dminus[222] = 18'b111111110_000011100;
		Dminus[223] = 18'b111111110_000011111;
		Dminus[224] = 18'b111111110_000100001;
		Dminus[225] = 18'b111111110_000100100;
		Dminus[226] = 18'b111111110_000100111;
		Dminus[227] = 18'b111111110_000101010;
		Dminus[228] = 18'b111111110_000101101;
		Dminus[229] = 18'b111111110_000101111;
		Dminus[230] = 18'b111111110_000110010;
		Dminus[231] = 18'b111111110_000110101;
		Dminus[232] = 18'b111111110_000111000;
		Dminus[233] = 18'b111111110_000111010;
		Dminus[234] = 18'b111111110_000111101;
		Dminus[235] = 18'b111111110_001000000;
		Dminus[236] = 18'b111111110_001000010;
		Dminus[237] = 18'b111111110_001000101;
		Dminus[238] = 18'b111111110_001001000;
		Dminus[239] = 18'b111111110_001001010;
		Dminus[240] = 18'b111111110_001001101;
		Dminus[241] = 18'b111111110_001001111;
		Dminus[242] = 18'b111111110_001010010;
		Dminus[243] = 18'b111111110_001010101;
		Dminus[244] = 18'b111111110_001010111;
		Dminus[245] = 18'b111111110_001011010;
		Dminus[246] = 18'b111111110_001011100;
		Dminus[247] = 18'b111111110_001011111;
		Dminus[248] = 18'b111111110_001100001;
		Dminus[249] = 18'b111111110_001100100;
		Dminus[250] = 18'b111111110_001100110;
		Dminus[251] = 18'b111111110_001101001;
		Dminus[252] = 18'b111111110_001101011;
		Dminus[253] = 18'b111111110_001101110;
		Dminus[254] = 18'b111111110_001110000;
		Dminus[255] = 18'b111111110_001110011;
		Dminus[256] = 18'b111111110_001110101;
		Dminus[257] = 18'b111111110_001110111;
		Dminus[258] = 18'b111111110_001111010;
		Dminus[259] = 18'b111111110_001111100;
		Dminus[260] = 18'b111111110_001111111;
		Dminus[261] = 18'b111111110_010000001;
		Dminus[262] = 18'b111111110_010000011;
		Dminus[263] = 18'b111111110_010000110;
		Dminus[264] = 18'b111111110_010001000;
		Dminus[265] = 18'b111111110_010001010;
		Dminus[266] = 18'b111111110_010001101;
		Dminus[267] = 18'b111111110_010001111;
		Dminus[268] = 18'b111111110_010010001;
		Dminus[269] = 18'b111111110_010010011;
		Dminus[270] = 18'b111111110_010010110;
		Dminus[271] = 18'b111111110_010011000;
		Dminus[272] = 18'b111111110_010011010;
		Dminus[273] = 18'b111111110_010011100;
		Dminus[274] = 18'b111111110_010011111;
		Dminus[275] = 18'b111111110_010100001;
		Dminus[276] = 18'b111111110_010100011;
		Dminus[277] = 18'b111111110_010100101;
		Dminus[278] = 18'b111111110_010101000;
		Dminus[279] = 18'b111111110_010101010;
		Dminus[280] = 18'b111111110_010101100;
		Dminus[281] = 18'b111111110_010101110;
		Dminus[282] = 18'b111111110_010110000;
		Dminus[283] = 18'b111111110_010110010;
		Dminus[284] = 18'b111111110_010110100;
		Dminus[285] = 18'b111111110_010110111;
		Dminus[286] = 18'b111111110_010111001;
		Dminus[287] = 18'b111111110_010111011;
		Dminus[288] = 18'b111111110_010111101;
		Dminus[289] = 18'b111111110_010111111;
		Dminus[290] = 18'b111111110_011000001;
		Dminus[291] = 18'b111111110_011000011;
		Dminus[292] = 18'b111111110_011000101;
		Dminus[293] = 18'b111111110_011000111;
		Dminus[294] = 18'b111111110_011001001;
		Dminus[295] = 18'b111111110_011001011;
		Dminus[296] = 18'b111111110_011001101;
		Dminus[297] = 18'b111111110_011001111;
		Dminus[298] = 18'b111111110_011010001;
		Dminus[299] = 18'b111111110_011010011;
		Dminus[300] = 18'b111111110_011010101;
		Dminus[301] = 18'b111111110_011010111;
		Dminus[302] = 18'b111111110_011011001;
		Dminus[303] = 18'b111111110_011011011;
		Dminus[304] = 18'b111111110_011011101;
		Dminus[305] = 18'b111111110_011011111;
		Dminus[306] = 18'b111111110_011100001;
		Dminus[307] = 18'b111111110_011100011;
		Dminus[308] = 18'b111111110_011100101;
		Dminus[309] = 18'b111111110_011100111;
		Dminus[310] = 18'b111111110_011101001;
		Dminus[311] = 18'b111111110_011101011;
		Dminus[312] = 18'b111111110_011101101;
		Dminus[313] = 18'b111111110_011101111;
		Dminus[314] = 18'b111111110_011110001;
		Dminus[315] = 18'b111111110_011110011;
		Dminus[316] = 18'b111111110_011110100;
		Dminus[317] = 18'b111111110_011110110;
		Dminus[318] = 18'b111111110_011111000;
		Dminus[319] = 18'b111111110_011111010;
		Dminus[320] = 18'b111111110_011111100;
		Dminus[321] = 18'b111111110_011111110;
		Dminus[322] = 18'b111111110_100000000;
		Dminus[323] = 18'b111111110_100000001;
		Dminus[324] = 18'b111111110_100000011;
		Dminus[325] = 18'b111111110_100000101;
		Dminus[326] = 18'b111111110_100000111;
		Dminus[327] = 18'b111111110_100001001;
		Dminus[328] = 18'b111111110_100001010;
		Dminus[329] = 18'b111111110_100001100;
		Dminus[330] = 18'b111111110_100001110;
		Dminus[331] = 18'b111111110_100010000;
		Dminus[332] = 18'b111111110_100010001;
		Dminus[333] = 18'b111111110_100010011;
		Dminus[334] = 18'b111111110_100010101;
		Dminus[335] = 18'b111111110_100010111;
		Dminus[336] = 18'b111111110_100011000;
		Dminus[337] = 18'b111111110_100011010;
		Dminus[338] = 18'b111111110_100011100;
		Dminus[339] = 18'b111111110_100011110;
		Dminus[340] = 18'b111111110_100011111;
		Dminus[341] = 18'b111111110_100100001;
		Dminus[342] = 18'b111111110_100100011;
		Dminus[343] = 18'b111111110_100100100;
		Dminus[344] = 18'b111111110_100100110;
		Dminus[345] = 18'b111111110_100101000;
		Dminus[346] = 18'b111111110_100101010;
		Dminus[347] = 18'b111111110_100101011;
		Dminus[348] = 18'b111111110_100101101;
		Dminus[349] = 18'b111111110_100101111;
		Dminus[350] = 18'b111111110_100110000;
		Dminus[351] = 18'b111111110_100110010;
		Dminus[352] = 18'b111111110_100110011;
		Dminus[353] = 18'b111111110_100110101;
		Dminus[354] = 18'b111111110_100110111;
		Dminus[355] = 18'b111111110_100111000;
		Dminus[356] = 18'b111111110_100111010;
		Dminus[357] = 18'b111111110_100111100;
		Dminus[358] = 18'b111111110_100111101;
		Dminus[359] = 18'b111111110_100111111;
		Dminus[360] = 18'b111111110_101000000;
		Dminus[361] = 18'b111111110_101000010;
		Dminus[362] = 18'b111111110_101000100;
		Dminus[363] = 18'b111111110_101000101;
		Dminus[364] = 18'b111111110_101000111;
		Dminus[365] = 18'b111111110_101001000;
		Dminus[366] = 18'b111111110_101001010;
		Dminus[367] = 18'b111111110_101001011;
		Dminus[368] = 18'b111111110_101001101;
		Dminus[369] = 18'b111111110_101001111;
		Dminus[370] = 18'b111111110_101010000;
		Dminus[371] = 18'b111111110_101010010;
		Dminus[372] = 18'b111111110_101010011;
		Dminus[373] = 18'b111111110_101010101;
		Dminus[374] = 18'b111111110_101010110;
		Dminus[375] = 18'b111111110_101011000;
		Dminus[376] = 18'b111111110_101011001;
		Dminus[377] = 18'b111111110_101011011;
		Dminus[378] = 18'b111111110_101011100;
		Dminus[379] = 18'b111111110_101011110;
		Dminus[380] = 18'b111111110_101011111;
		Dminus[381] = 18'b111111110_101100001;
		Dminus[382] = 18'b111111110_101100010;
		Dminus[383] = 18'b111111110_101100100;
		Dminus[384] = 18'b111111110_101100101;
		Dminus[385] = 18'b111111110_101100111;
		Dminus[386] = 18'b111111110_101101000;
		Dminus[387] = 18'b111111110_101101001;
		Dminus[388] = 18'b111111110_101101011;
		Dminus[389] = 18'b111111110_101101100;
		Dminus[390] = 18'b111111110_101101110;
		Dminus[391] = 18'b111111110_101101111;
		Dminus[392] = 18'b111111110_101110001;
		Dminus[393] = 18'b111111110_101110010;
		Dminus[394] = 18'b111111110_101110011;
		Dminus[395] = 18'b111111110_101110101;
		Dminus[396] = 18'b111111110_101110110;
		Dminus[397] = 18'b111111110_101111000;
		Dminus[398] = 18'b111111110_101111001;
		Dminus[399] = 18'b111111110_101111011;
		Dminus[400] = 18'b111111110_101111100;
		Dminus[401] = 18'b111111110_101111101;
		Dminus[402] = 18'b111111110_101111111;
		Dminus[403] = 18'b111111110_110000000;
		Dminus[404] = 18'b111111110_110000001;
		Dminus[405] = 18'b111111110_110000011;
		Dminus[406] = 18'b111111110_110000100;
		Dminus[407] = 18'b111111110_110000110;
		Dminus[408] = 18'b111111110_110000111;
		Dminus[409] = 18'b111111110_110001000;
		Dminus[410] = 18'b111111110_110001010;
		Dminus[411] = 18'b111111110_110001011;
		Dminus[412] = 18'b111111110_110001100;
		Dminus[413] = 18'b111111110_110001110;
		Dminus[414] = 18'b111111110_110001111;
		Dminus[415] = 18'b111111110_110010000;
		Dminus[416] = 18'b111111110_110010010;
		Dminus[417] = 18'b111111110_110010011;
		Dminus[418] = 18'b111111110_110010100;
		Dminus[419] = 18'b111111110_110010110;
		Dminus[420] = 18'b111111110_110010111;
		Dminus[421] = 18'b111111110_110011000;
		Dminus[422] = 18'b111111110_110011001;
		Dminus[423] = 18'b111111110_110011011;
		Dminus[424] = 18'b111111110_110011100;
		Dminus[425] = 18'b111111110_110011101;
		Dminus[426] = 18'b111111110_110011111;
		Dminus[427] = 18'b111111110_110100000;
		Dminus[428] = 18'b111111110_110100001;
		Dminus[429] = 18'b111111110_110100010;
		Dminus[430] = 18'b111111110_110100100;
		Dminus[431] = 18'b111111110_110100101;
		Dminus[432] = 18'b111111110_110100110;
		Dminus[433] = 18'b111111110_110101000;
		Dminus[434] = 18'b111111110_110101001;
		Dminus[435] = 18'b111111110_110101010;
		Dminus[436] = 18'b111111110_110101011;
		Dminus[437] = 18'b111111110_110101101;
		Dminus[438] = 18'b111111110_110101110;
		Dminus[439] = 18'b111111110_110101111;
		Dminus[440] = 18'b111111110_110110000;
		Dminus[441] = 18'b111111110_110110001;
		Dminus[442] = 18'b111111110_110110011;
		Dminus[443] = 18'b111111110_110110100;
		Dminus[444] = 18'b111111110_110110101;
		Dminus[445] = 18'b111111110_110110110;
		Dminus[446] = 18'b111111110_110111000;
		Dminus[447] = 18'b111111110_110111001;
		Dminus[448] = 18'b111111110_110111010;
		Dminus[449] = 18'b111111110_110111011;
		Dminus[450] = 18'b111111110_110111100;
		Dminus[451] = 18'b111111110_110111110;
		Dminus[452] = 18'b111111110_110111111;
		Dminus[453] = 18'b111111110_111000000;
		Dminus[454] = 18'b111111110_111000001;
		Dminus[455] = 18'b111111110_111000010;
		Dminus[456] = 18'b111111110_111000011;
		Dminus[457] = 18'b111111110_111000101;
		Dminus[458] = 18'b111111110_111000110;
		Dminus[459] = 18'b111111110_111000111;
		Dminus[460] = 18'b111111110_111001000;
		Dminus[461] = 18'b111111110_111001001;
		Dminus[462] = 18'b111111110_111001010;
		Dminus[463] = 18'b111111110_111001100;
		Dminus[464] = 18'b111111110_111001101;
		Dminus[465] = 18'b111111110_111001110;
		Dminus[466] = 18'b111111110_111001111;
		Dminus[467] = 18'b111111110_111010000;
		Dminus[468] = 18'b111111110_111010001;
		Dminus[469] = 18'b111111110_111010010;
		Dminus[470] = 18'b111111110_111010011;
		Dminus[471] = 18'b111111110_111010101;
		Dminus[472] = 18'b111111110_111010110;
		Dminus[473] = 18'b111111110_111010111;
		Dminus[474] = 18'b111111110_111011000;
		Dminus[475] = 18'b111111110_111011001;
		Dminus[476] = 18'b111111110_111011010;
		Dminus[477] = 18'b111111110_111011011;
		Dminus[478] = 18'b111111110_111011100;
		Dminus[479] = 18'b111111110_111011101;
		Dminus[480] = 18'b111111110_111011111;
		Dminus[481] = 18'b111111110_111100000;
		Dminus[482] = 18'b111111110_111100001;
		Dminus[483] = 18'b111111110_111100010;
		Dminus[484] = 18'b111111110_111100011;
		Dminus[485] = 18'b111111110_111100100;
		Dminus[486] = 18'b111111110_111100101;
		Dminus[487] = 18'b111111110_111100110;
		Dminus[488] = 18'b111111110_111100111;
		Dminus[489] = 18'b111111110_111101000;
		Dminus[490] = 18'b111111110_111101001;
		Dminus[491] = 18'b111111110_111101010;
		Dminus[492] = 18'b111111110_111101011;
		Dminus[493] = 18'b111111110_111101100;
		Dminus[494] = 18'b111111110_111101110;
		Dminus[495] = 18'b111111110_111101111;
		Dminus[496] = 18'b111111110_111110000;
		Dminus[497] = 18'b111111110_111110001;
		Dminus[498] = 18'b111111110_111110010;
		Dminus[499] = 18'b111111110_111110011;
		Dminus[500] = 18'b111111110_111110100;
		Dminus[501] = 18'b111111110_111110101;
		Dminus[502] = 18'b111111110_111110110;
		Dminus[503] = 18'b111111110_111110111;
		Dminus[504] = 18'b111111110_111111000;
		Dminus[505] = 18'b111111110_111111001;
		Dminus[506] = 18'b111111110_111111010;
		Dminus[507] = 18'b111111110_111111011;
		Dminus[508] = 18'b111111110_111111100;
		Dminus[509] = 18'b111111110_111111101;
		Dminus[510] = 18'b111111110_111111110;
		Dminus[511] = 18'b111111110_111111111;
		Dminus[512] = 18'b111111111_000000000;
		Dminus[513] = 18'b111111111_000000001;
		Dminus[514] = 18'b111111111_000000010;
		Dminus[515] = 18'b111111111_000000011;
		Dminus[516] = 18'b111111111_000000100;
		Dminus[517] = 18'b111111111_000000101;
		Dminus[518] = 18'b111111111_000000110;
		Dminus[519] = 18'b111111111_000000111;
		Dminus[520] = 18'b111111111_000001000;
		Dminus[521] = 18'b111111111_000001001;
		Dminus[522] = 18'b111111111_000001010;
		Dminus[523] = 18'b111111111_000001011;
		Dminus[524] = 18'b111111111_000001100;
		Dminus[525] = 18'b111111111_000001101;
		Dminus[526] = 18'b111111111_000001110;
		Dminus[527] = 18'b111111111_000001111;
		Dminus[528] = 18'b111111111_000010000;
		Dminus[529] = 18'b111111111_000010001;
		Dminus[530] = 18'b111111111_000010010;
		Dminus[531] = 18'b111111111_000010011;
		Dminus[532] = 18'b111111111_000010011;
		Dminus[533] = 18'b111111111_000010100;
		Dminus[534] = 18'b111111111_000010101;
		Dminus[535] = 18'b111111111_000010110;
		Dminus[536] = 18'b111111111_000010111;
		Dminus[537] = 18'b111111111_000011000;
		Dminus[538] = 18'b111111111_000011001;
		Dminus[539] = 18'b111111111_000011010;
		Dminus[540] = 18'b111111111_000011011;
		Dminus[541] = 18'b111111111_000011100;
		Dminus[542] = 18'b111111111_000011101;
		Dminus[543] = 18'b111111111_000011110;
		Dminus[544] = 18'b111111111_000011111;
		Dminus[545] = 18'b111111111_000100000;
		Dminus[546] = 18'b111111111_000100001;
		Dminus[547] = 18'b111111111_000100001;
		Dminus[548] = 18'b111111111_000100010;
		Dminus[549] = 18'b111111111_000100011;
		Dminus[550] = 18'b111111111_000100100;
		Dminus[551] = 18'b111111111_000100101;
		Dminus[552] = 18'b111111111_000100110;
		Dminus[553] = 18'b111111111_000100111;
		Dminus[554] = 18'b111111111_000101000;
		Dminus[555] = 18'b111111111_000101001;
		Dminus[556] = 18'b111111111_000101010;
		Dminus[557] = 18'b111111111_000101010;
		Dminus[558] = 18'b111111111_000101011;
		Dminus[559] = 18'b111111111_000101100;
		Dminus[560] = 18'b111111111_000101101;
		Dminus[561] = 18'b111111111_000101110;
		Dminus[562] = 18'b111111111_000101111;
		Dminus[563] = 18'b111111111_000110000;
		Dminus[564] = 18'b111111111_000110001;
		Dminus[565] = 18'b111111111_000110001;
		Dminus[566] = 18'b111111111_000110010;
		Dminus[567] = 18'b111111111_000110011;
		Dminus[568] = 18'b111111111_000110100;
		Dminus[569] = 18'b111111111_000110101;
		Dminus[570] = 18'b111111111_000110110;
		Dminus[571] = 18'b111111111_000110111;
		Dminus[572] = 18'b111111111_000110111;
		Dminus[573] = 18'b111111111_000111000;
		Dminus[574] = 18'b111111111_000111001;
		Dminus[575] = 18'b111111111_000111010;
		Dminus[576] = 18'b111111111_000111011;
		Dminus[577] = 18'b111111111_000111100;
		Dminus[578] = 18'b111111111_000111101;
		Dminus[579] = 18'b111111111_000111101;
		Dminus[580] = 18'b111111111_000111110;
		Dminus[581] = 18'b111111111_000111111;
		Dminus[582] = 18'b111111111_001000000;
		Dminus[583] = 18'b111111111_001000001;
		Dminus[584] = 18'b111111111_001000010;
		Dminus[585] = 18'b111111111_001000010;
		Dminus[586] = 18'b111111111_001000011;
		Dminus[587] = 18'b111111111_001000100;
		Dminus[588] = 18'b111111111_001000101;
		Dminus[589] = 18'b111111111_001000110;
		Dminus[590] = 18'b111111111_001000111;
		Dminus[591] = 18'b111111111_001000111;
		Dminus[592] = 18'b111111111_001001000;
		Dminus[593] = 18'b111111111_001001001;
		Dminus[594] = 18'b111111111_001001010;
		Dminus[595] = 18'b111111111_001001011;
		Dminus[596] = 18'b111111111_001001011;
		Dminus[597] = 18'b111111111_001001100;
		Dminus[598] = 18'b111111111_001001101;
		Dminus[599] = 18'b111111111_001001110;
		Dminus[600] = 18'b111111111_001001111;
		Dminus[601] = 18'b111111111_001001111;
		Dminus[602] = 18'b111111111_001010000;
		Dminus[603] = 18'b111111111_001010001;
		Dminus[604] = 18'b111111111_001010010;
		Dminus[605] = 18'b111111111_001010011;
		Dminus[606] = 18'b111111111_001010011;
		Dminus[607] = 18'b111111111_001010100;
		Dminus[608] = 18'b111111111_001010101;
		Dminus[609] = 18'b111111111_001010110;
		Dminus[610] = 18'b111111111_001010111;
		Dminus[611] = 18'b111111111_001010111;
		Dminus[612] = 18'b111111111_001011000;
		Dminus[613] = 18'b111111111_001011001;
		Dminus[614] = 18'b111111111_001011010;
		Dminus[615] = 18'b111111111_001011010;
		Dminus[616] = 18'b111111111_001011011;
		Dminus[617] = 18'b111111111_001011100;
		Dminus[618] = 18'b111111111_001011101;
		Dminus[619] = 18'b111111111_001011101;
		Dminus[620] = 18'b111111111_001011110;
		Dminus[621] = 18'b111111111_001011111;
		Dminus[622] = 18'b111111111_001100000;
		Dminus[623] = 18'b111111111_001100000;
		Dminus[624] = 18'b111111111_001100001;
		Dminus[625] = 18'b111111111_001100010;
		Dminus[626] = 18'b111111111_001100011;
		Dminus[627] = 18'b111111111_001100011;
		Dminus[628] = 18'b111111111_001100100;
		Dminus[629] = 18'b111111111_001100101;
		Dminus[630] = 18'b111111111_001100110;
		Dminus[631] = 18'b111111111_001100110;
		Dminus[632] = 18'b111111111_001100111;
		Dminus[633] = 18'b111111111_001101000;
		Dminus[634] = 18'b111111111_001101001;
		Dminus[635] = 18'b111111111_001101001;
		Dminus[636] = 18'b111111111_001101010;
		Dminus[637] = 18'b111111111_001101011;
		Dminus[638] = 18'b111111111_001101100;
		Dminus[639] = 18'b111111111_001101100;
		Dminus[640] = 18'b111111111_001101101;
		Dminus[641] = 18'b111111111_001101110;
		Dminus[642] = 18'b111111111_001101111;
		Dminus[643] = 18'b111111111_001101111;
		Dminus[644] = 18'b111111111_001110000;
		Dminus[645] = 18'b111111111_001110001;
		Dminus[646] = 18'b111111111_001110001;
		Dminus[647] = 18'b111111111_001110010;
		Dminus[648] = 18'b111111111_001110011;
		Dminus[649] = 18'b111111111_001110100;
		Dminus[650] = 18'b111111111_001110100;
		Dminus[651] = 18'b111111111_001110101;
		Dminus[652] = 18'b111111111_001110110;
		Dminus[653] = 18'b111111111_001110110;
		Dminus[654] = 18'b111111111_001110111;
		Dminus[655] = 18'b111111111_001111000;
		Dminus[656] = 18'b111111111_001111000;
		Dminus[657] = 18'b111111111_001111001;
		Dminus[658] = 18'b111111111_001111010;
		Dminus[659] = 18'b111111111_001111011;
		Dminus[660] = 18'b111111111_001111011;
		Dminus[661] = 18'b111111111_001111100;
		Dminus[662] = 18'b111111111_001111101;
		Dminus[663] = 18'b111111111_001111101;
		Dminus[664] = 18'b111111111_001111110;
		Dminus[665] = 18'b111111111_001111111;
		Dminus[666] = 18'b111111111_001111111;
		Dminus[667] = 18'b111111111_010000000;
		Dminus[668] = 18'b111111111_010000001;
		Dminus[669] = 18'b111111111_010000001;
		Dminus[670] = 18'b111111111_010000010;
		Dminus[671] = 18'b111111111_010000011;
		Dminus[672] = 18'b111111111_010000011;
		Dminus[673] = 18'b111111111_010000100;
		Dminus[674] = 18'b111111111_010000101;
		Dminus[675] = 18'b111111111_010000101;
		Dminus[676] = 18'b111111111_010000110;
		Dminus[677] = 18'b111111111_010000111;
		Dminus[678] = 18'b111111111_010000111;
		Dminus[679] = 18'b111111111_010001000;
		Dminus[680] = 18'b111111111_010001001;
		Dminus[681] = 18'b111111111_010001001;
		Dminus[682] = 18'b111111111_010001010;
		Dminus[683] = 18'b111111111_010001011;
		Dminus[684] = 18'b111111111_010001011;
		Dminus[685] = 18'b111111111_010001100;
		Dminus[686] = 18'b111111111_010001101;
		Dminus[687] = 18'b111111111_010001101;
		Dminus[688] = 18'b111111111_010001110;
		Dminus[689] = 18'b111111111_010001111;
		Dminus[690] = 18'b111111111_010001111;
		Dminus[691] = 18'b111111111_010010000;
		Dminus[692] = 18'b111111111_010010001;
		Dminus[693] = 18'b111111111_010010001;
		Dminus[694] = 18'b111111111_010010010;
		Dminus[695] = 18'b111111111_010010011;
		Dminus[696] = 18'b111111111_010010011;
		Dminus[697] = 18'b111111111_010010100;
		Dminus[698] = 18'b111111111_010010100;
		Dminus[699] = 18'b111111111_010010101;
		Dminus[700] = 18'b111111111_010010110;
		Dminus[701] = 18'b111111111_010010110;
		Dminus[702] = 18'b111111111_010010111;
		Dminus[703] = 18'b111111111_010011000;
		Dminus[704] = 18'b111111111_010011000;
		Dminus[705] = 18'b111111111_010011001;
		Dminus[706] = 18'b111111111_010011010;
		Dminus[707] = 18'b111111111_010011010;
		Dminus[708] = 18'b111111111_010011011;
		Dminus[709] = 18'b111111111_010011011;
		Dminus[710] = 18'b111111111_010011100;
		Dminus[711] = 18'b111111111_010011101;
		Dminus[712] = 18'b111111111_010011101;
		Dminus[713] = 18'b111111111_010011110;
		Dminus[714] = 18'b111111111_010011110;
		Dminus[715] = 18'b111111111_010011111;
		Dminus[716] = 18'b111111111_010100000;
		Dminus[717] = 18'b111111111_010100000;
		Dminus[718] = 18'b111111111_010100001;
		Dminus[719] = 18'b111111111_010100010;
		Dminus[720] = 18'b111111111_010100010;
		Dminus[721] = 18'b111111111_010100011;
		Dminus[722] = 18'b111111111_010100011;
		Dminus[723] = 18'b111111111_010100100;
		Dminus[724] = 18'b111111111_010100101;
		Dminus[725] = 18'b111111111_010100101;
		Dminus[726] = 18'b111111111_010100110;
		Dminus[727] = 18'b111111111_010100110;
		Dminus[728] = 18'b111111111_010100111;
		Dminus[729] = 18'b111111111_010101000;
		Dminus[730] = 18'b111111111_010101000;
		Dminus[731] = 18'b111111111_010101001;
		Dminus[732] = 18'b111111111_010101001;
		Dminus[733] = 18'b111111111_010101010;
		Dminus[734] = 18'b111111111_010101010;
		Dminus[735] = 18'b111111111_010101011;
		Dminus[736] = 18'b111111111_010101100;
		Dminus[737] = 18'b111111111_010101100;
		Dminus[738] = 18'b111111111_010101101;
		Dminus[739] = 18'b111111111_010101101;
		Dminus[740] = 18'b111111111_010101110;
		Dminus[741] = 18'b111111111_010101111;
		Dminus[742] = 18'b111111111_010101111;
		Dminus[743] = 18'b111111111_010110000;
		Dminus[744] = 18'b111111111_010110000;
		Dminus[745] = 18'b111111111_010110001;
		Dminus[746] = 18'b111111111_010110001;
		Dminus[747] = 18'b111111111_010110010;
		Dminus[748] = 18'b111111111_010110011;
		Dminus[749] = 18'b111111111_010110011;
		Dminus[750] = 18'b111111111_010110100;
		Dminus[751] = 18'b111111111_010110100;
		Dminus[752] = 18'b111111111_010110101;
		Dminus[753] = 18'b111111111_010110101;
		Dminus[754] = 18'b111111111_010110110;
		Dminus[755] = 18'b111111111_010110111;
		Dminus[756] = 18'b111111111_010110111;
		Dminus[757] = 18'b111111111_010111000;
		Dminus[758] = 18'b111111111_010111000;
		Dminus[759] = 18'b111111111_010111001;
		Dminus[760] = 18'b111111111_010111001;
		Dminus[761] = 18'b111111111_010111010;
		Dminus[762] = 18'b111111111_010111010;
		Dminus[763] = 18'b111111111_010111011;
		Dminus[764] = 18'b111111111_010111100;
		Dminus[765] = 18'b111111111_010111100;
		Dminus[766] = 18'b111111111_010111101;
		Dminus[767] = 18'b111111111_010111101;
		Dminus[768] = 18'b111111111_010111110;
		Dminus[769] = 18'b111111111_010111110;
		Dminus[770] = 18'b111111111_010111111;
		Dminus[771] = 18'b111111111_010111111;
		Dminus[772] = 18'b111111111_011000000;
		Dminus[773] = 18'b111111111_011000000;
		Dminus[774] = 18'b111111111_011000001;
		Dminus[775] = 18'b111111111_011000010;
		Dminus[776] = 18'b111111111_011000010;
		Dminus[777] = 18'b111111111_011000011;
		Dminus[778] = 18'b111111111_011000011;
		Dminus[779] = 18'b111111111_011000100;
		Dminus[780] = 18'b111111111_011000100;
		Dminus[781] = 18'b111111111_011000101;
		Dminus[782] = 18'b111111111_011000101;
		Dminus[783] = 18'b111111111_011000110;
		Dminus[784] = 18'b111111111_011000110;
		Dminus[785] = 18'b111111111_011000111;
		Dminus[786] = 18'b111111111_011000111;
		Dminus[787] = 18'b111111111_011001000;
		Dminus[788] = 18'b111111111_011001000;
		Dminus[789] = 18'b111111111_011001001;
		Dminus[790] = 18'b111111111_011001010;
		Dminus[791] = 18'b111111111_011001010;
		Dminus[792] = 18'b111111111_011001011;
		Dminus[793] = 18'b111111111_011001011;
		Dminus[794] = 18'b111111111_011001100;
		Dminus[795] = 18'b111111111_011001100;
		Dminus[796] = 18'b111111111_011001101;
		Dminus[797] = 18'b111111111_011001101;
		Dminus[798] = 18'b111111111_011001110;
		Dminus[799] = 18'b111111111_011001110;
		Dminus[800] = 18'b111111111_011001111;
		Dminus[801] = 18'b111111111_011001111;
		Dminus[802] = 18'b111111111_011010000;
		Dminus[803] = 18'b111111111_011010000;
		Dminus[804] = 18'b111111111_011010001;
		Dminus[805] = 18'b111111111_011010001;
		Dminus[806] = 18'b111111111_011010010;
		Dminus[807] = 18'b111111111_011010010;
		Dminus[808] = 18'b111111111_011010011;
		Dminus[809] = 18'b111111111_011010011;
		Dminus[810] = 18'b111111111_011010100;
		Dminus[811] = 18'b111111111_011010100;
		Dminus[812] = 18'b111111111_011010101;
		Dminus[813] = 18'b111111111_011010101;
		Dminus[814] = 18'b111111111_011010110;
		Dminus[815] = 18'b111111111_011010110;
		Dminus[816] = 18'b111111111_011010111;
		Dminus[817] = 18'b111111111_011010111;
		Dminus[818] = 18'b111111111_011011000;
		Dminus[819] = 18'b111111111_011011000;
		Dminus[820] = 18'b111111111_011011001;
		Dminus[821] = 18'b111111111_011011001;
		Dminus[822] = 18'b111111111_011011010;
		Dminus[823] = 18'b111111111_011011010;
		Dminus[824] = 18'b111111111_011011011;
		Dminus[825] = 18'b111111111_011011011;
		Dminus[826] = 18'b111111111_011011100;
		Dminus[827] = 18'b111111111_011011100;
		Dminus[828] = 18'b111111111_011011101;
		Dminus[829] = 18'b111111111_011011101;
		Dminus[830] = 18'b111111111_011011110;
		Dminus[831] = 18'b111111111_011011110;
		Dminus[832] = 18'b111111111_011011111;
		Dminus[833] = 18'b111111111_011011111;
		Dminus[834] = 18'b111111111_011011111;
		Dminus[835] = 18'b111111111_011100000;
		Dminus[836] = 18'b111111111_011100000;
		Dminus[837] = 18'b111111111_011100001;
		Dminus[838] = 18'b111111111_011100001;
		Dminus[839] = 18'b111111111_011100010;
		Dminus[840] = 18'b111111111_011100010;
		Dminus[841] = 18'b111111111_011100011;
		Dminus[842] = 18'b111111111_011100011;
		Dminus[843] = 18'b111111111_011100100;
		Dminus[844] = 18'b111111111_011100100;
		Dminus[845] = 18'b111111111_011100101;
		Dminus[846] = 18'b111111111_011100101;
		Dminus[847] = 18'b111111111_011100110;
		Dminus[848] = 18'b111111111_011100110;
		Dminus[849] = 18'b111111111_011100111;
		Dminus[850] = 18'b111111111_011100111;
		Dminus[851] = 18'b111111111_011100111;
		Dminus[852] = 18'b111111111_011101000;
		Dminus[853] = 18'b111111111_011101000;
		Dminus[854] = 18'b111111111_011101001;
		Dminus[855] = 18'b111111111_011101001;
		Dminus[856] = 18'b111111111_011101010;
		Dminus[857] = 18'b111111111_011101010;
		Dminus[858] = 18'b111111111_011101011;
		Dminus[859] = 18'b111111111_011101011;
		Dminus[860] = 18'b111111111_011101100;
		Dminus[861] = 18'b111111111_011101100;
		Dminus[862] = 18'b111111111_011101101;
		Dminus[863] = 18'b111111111_011101101;
		Dminus[864] = 18'b111111111_011101101;
		Dminus[865] = 18'b111111111_011101110;
		Dminus[866] = 18'b111111111_011101110;
		Dminus[867] = 18'b111111111_011101111;
		Dminus[868] = 18'b111111111_011101111;
		Dminus[869] = 18'b111111111_011110000;
		Dminus[870] = 18'b111111111_011110000;
		Dminus[871] = 18'b111111111_011110001;
		Dminus[872] = 18'b111111111_011110001;
		Dminus[873] = 18'b111111111_011110001;
		Dminus[874] = 18'b111111111_011110010;
		Dminus[875] = 18'b111111111_011110010;
		Dminus[876] = 18'b111111111_011110011;
		Dminus[877] = 18'b111111111_011110011;
		Dminus[878] = 18'b111111111_011110100;
		Dminus[879] = 18'b111111111_011110100;
		Dminus[880] = 18'b111111111_011110101;
		Dminus[881] = 18'b111111111_011110101;
		Dminus[882] = 18'b111111111_011110101;
		Dminus[883] = 18'b111111111_011110110;
		Dminus[884] = 18'b111111111_011110110;
		Dminus[885] = 18'b111111111_011110111;
		Dminus[886] = 18'b111111111_011110111;
		Dminus[887] = 18'b111111111_011111000;
		Dminus[888] = 18'b111111111_011111000;
		Dminus[889] = 18'b111111111_011111000;
		Dminus[890] = 18'b111111111_011111001;
		Dminus[891] = 18'b111111111_011111001;
		Dminus[892] = 18'b111111111_011111010;
		Dminus[893] = 18'b111111111_011111010;
		Dminus[894] = 18'b111111111_011111011;
		Dminus[895] = 18'b111111111_011111011;
		Dminus[896] = 18'b111111111_011111011;
		Dminus[897] = 18'b111111111_011111100;
		Dminus[898] = 18'b111111111_011111100;
		Dminus[899] = 18'b111111111_011111101;
		Dminus[900] = 18'b111111111_011111101;
		Dminus[901] = 18'b111111111_011111101;
		Dminus[902] = 18'b111111111_011111110;
		Dminus[903] = 18'b111111111_011111110;
		Dminus[904] = 18'b111111111_011111111;
		Dminus[905] = 18'b111111111_011111111;
		Dminus[906] = 18'b111111111_100000000;
		Dminus[907] = 18'b111111111_100000000;
		Dminus[908] = 18'b111111111_100000000;
		Dminus[909] = 18'b111111111_100000001;
		Dminus[910] = 18'b111111111_100000001;
		Dminus[911] = 18'b111111111_100000010;
		Dminus[912] = 18'b111111111_100000010;
		Dminus[913] = 18'b111111111_100000010;
		Dminus[914] = 18'b111111111_100000011;
		Dminus[915] = 18'b111111111_100000011;
		Dminus[916] = 18'b111111111_100000100;
		Dminus[917] = 18'b111111111_100000100;
		Dminus[918] = 18'b111111111_100000100;
		Dminus[919] = 18'b111111111_100000101;
		Dminus[920] = 18'b111111111_100000101;
		Dminus[921] = 18'b111111111_100000110;
		Dminus[922] = 18'b111111111_100000110;
		Dminus[923] = 18'b111111111_100000111;
		Dminus[924] = 18'b111111111_100000111;
		Dminus[925] = 18'b111111111_100000111;
		Dminus[926] = 18'b111111111_100001000;
		Dminus[927] = 18'b111111111_100001000;
		Dminus[928] = 18'b111111111_100001001;
		Dminus[929] = 18'b111111111_100001001;
		Dminus[930] = 18'b111111111_100001001;
		Dminus[931] = 18'b111111111_100001010;
		Dminus[932] = 18'b111111111_100001010;
		Dminus[933] = 18'b111111111_100001010;
		Dminus[934] = 18'b111111111_100001011;
		Dminus[935] = 18'b111111111_100001011;
		Dminus[936] = 18'b111111111_100001100;
		Dminus[937] = 18'b111111111_100001100;
		Dminus[938] = 18'b111111111_100001100;
		Dminus[939] = 18'b111111111_100001101;
		Dminus[940] = 18'b111111111_100001101;
		Dminus[941] = 18'b111111111_100001110;
		Dminus[942] = 18'b111111111_100001110;
		Dminus[943] = 18'b111111111_100001110;
		Dminus[944] = 18'b111111111_100001111;
		Dminus[945] = 18'b111111111_100001111;
		Dminus[946] = 18'b111111111_100010000;
		Dminus[947] = 18'b111111111_100010000;
		Dminus[948] = 18'b111111111_100010000;
		Dminus[949] = 18'b111111111_100010001;
		Dminus[950] = 18'b111111111_100010001;
		Dminus[951] = 18'b111111111_100010001;
		Dminus[952] = 18'b111111111_100010010;
		Dminus[953] = 18'b111111111_100010010;
		Dminus[954] = 18'b111111111_100010011;
		Dminus[955] = 18'b111111111_100010011;
		Dminus[956] = 18'b111111111_100010011;
		Dminus[957] = 18'b111111111_100010100;
		Dminus[958] = 18'b111111111_100010100;
		Dminus[959] = 18'b111111111_100010100;
		Dminus[960] = 18'b111111111_100010101;
		Dminus[961] = 18'b111111111_100010101;
		Dminus[962] = 18'b111111111_100010110;
		Dminus[963] = 18'b111111111_100010110;
		Dminus[964] = 18'b111111111_100010110;
		Dminus[965] = 18'b111111111_100010111;
		Dminus[966] = 18'b111111111_100010111;
		Dminus[967] = 18'b111111111_100010111;
		Dminus[968] = 18'b111111111_100011000;
		Dminus[969] = 18'b111111111_100011000;
		Dminus[970] = 18'b111111111_100011001;
		Dminus[971] = 18'b111111111_100011001;
		Dminus[972] = 18'b111111111_100011001;
		Dminus[973] = 18'b111111111_100011010;
		Dminus[974] = 18'b111111111_100011010;
		Dminus[975] = 18'b111111111_100011010;
		Dminus[976] = 18'b111111111_100011011;
		Dminus[977] = 18'b111111111_100011011;
		Dminus[978] = 18'b111111111_100011100;
		Dminus[979] = 18'b111111111_100011100;
		Dminus[980] = 18'b111111111_100011100;
		Dminus[981] = 18'b111111111_100011101;
		Dminus[982] = 18'b111111111_100011101;
		Dminus[983] = 18'b111111111_100011101;
		Dminus[984] = 18'b111111111_100011110;
		Dminus[985] = 18'b111111111_100011110;
		Dminus[986] = 18'b111111111_100011110;
		Dminus[987] = 18'b111111111_100011111;
		Dminus[988] = 18'b111111111_100011111;
		Dminus[989] = 18'b111111111_100011111;
		Dminus[990] = 18'b111111111_100100000;
		Dminus[991] = 18'b111111111_100100000;
		Dminus[992] = 18'b111111111_100100001;
		Dminus[993] = 18'b111111111_100100001;
		Dminus[994] = 18'b111111111_100100001;
		Dminus[995] = 18'b111111111_100100010;
		Dminus[996] = 18'b111111111_100100010;
		Dminus[997] = 18'b111111111_100100010;
		Dminus[998] = 18'b111111111_100100011;
		Dminus[999] = 18'b111111111_100100011;
		Dminus[1000] = 18'b111111111_100100011;
		Dminus[1001] = 18'b111111111_100100100;
		Dminus[1002] = 18'b111111111_100100100;
		Dminus[1003] = 18'b111111111_100100100;
		Dminus[1004] = 18'b111111111_100100101;
		Dminus[1005] = 18'b111111111_100100101;
		Dminus[1006] = 18'b111111111_100100101;
		Dminus[1007] = 18'b111111111_100100110;
		Dminus[1008] = 18'b111111111_100100110;
		Dminus[1009] = 18'b111111111_100100110;
		Dminus[1010] = 18'b111111111_100100111;
		Dminus[1011] = 18'b111111111_100100111;
		Dminus[1012] = 18'b111111111_100100111;
		Dminus[1013] = 18'b111111111_100101000;
		Dminus[1014] = 18'b111111111_100101000;
		Dminus[1015] = 18'b111111111_100101000;
		Dminus[1016] = 18'b111111111_100101001;
		Dminus[1017] = 18'b111111111_100101001;
		Dminus[1018] = 18'b111111111_100101001;
		Dminus[1019] = 18'b111111111_100101010;
		Dminus[1020] = 18'b111111111_100101010;
		Dminus[1021] = 18'b111111111_100101010;
		Dminus[1022] = 18'b111111111_100101011;
		Dminus[1023] = 18'b111111111_100101011;
		Dplus[1] = 18'b000000001_000000000;
		Dplus[2] = 18'b000000000_111111111;
		Dplus[3] = 18'b000000000_111111111;
		Dplus[4] = 18'b000000000_111111110;
		Dplus[5] = 18'b000000000_111111110;
		Dplus[6] = 18'b000000000_111111101;
		Dplus[7] = 18'b000000000_111111101;
		Dplus[8] = 18'b000000000_111111100;
		Dplus[9] = 18'b000000000_111111100;
		Dplus[10] = 18'b000000000_111111011;
		Dplus[11] = 18'b000000000_111111011;
		Dplus[12] = 18'b000000000_111111010;
		Dplus[13] = 18'b000000000_111111010;
		Dplus[14] = 18'b000000000_111111001;
		Dplus[15] = 18'b000000000_111111001;
		Dplus[16] = 18'b000000000_111111000;
		Dplus[17] = 18'b000000000_111111000;
		Dplus[18] = 18'b000000000_111110111;
		Dplus[19] = 18'b000000000_111110111;
		Dplus[20] = 18'b000000000_111110110;
		Dplus[21] = 18'b000000000_111110110;
		Dplus[22] = 18'b000000000_111110101;
		Dplus[23] = 18'b000000000_111110101;
		Dplus[24] = 18'b000000000_111110100;
		Dplus[25] = 18'b000000000_111110100;
		Dplus[26] = 18'b000000000_111110011;
		Dplus[27] = 18'b000000000_111110011;
		Dplus[28] = 18'b000000000_111110010;
		Dplus[29] = 18'b000000000_111110010;
		Dplus[30] = 18'b000000000_111110001;
		Dplus[31] = 18'b000000000_111110001;
		Dplus[32] = 18'b000000000_111110000;
		Dplus[33] = 18'b000000000_111110000;
		Dplus[34] = 18'b000000000_111101111;
		Dplus[35] = 18'b000000000_111101111;
		Dplus[36] = 18'b000000000_111101110;
		Dplus[37] = 18'b000000000_111101110;
		Dplus[38] = 18'b000000000_111101101;
		Dplus[39] = 18'b000000000_111101101;
		Dplus[40] = 18'b000000000_111101100;
		Dplus[41] = 18'b000000000_111101100;
		Dplus[42] = 18'b000000000_111101011;
		Dplus[43] = 18'b000000000_111101011;
		Dplus[44] = 18'b000000000_111101010;
		Dplus[45] = 18'b000000000_111101010;
		Dplus[46] = 18'b000000000_111101001;
		Dplus[47] = 18'b000000000_111101001;
		Dplus[48] = 18'b000000000_111101000;
		Dplus[49] = 18'b000000000_111101000;
		Dplus[50] = 18'b000000000_111100111;
		Dplus[51] = 18'b000000000_111100111;
		Dplus[52] = 18'b000000000_111100110;
		Dplus[53] = 18'b000000000_111100110;
		Dplus[54] = 18'b000000000_111100101;
		Dplus[55] = 18'b000000000_111100101;
		Dplus[56] = 18'b000000000_111100101;
		Dplus[57] = 18'b000000000_111100100;
		Dplus[58] = 18'b000000000_111100100;
		Dplus[59] = 18'b000000000_111100011;
		Dplus[60] = 18'b000000000_111100011;
		Dplus[61] = 18'b000000000_111100010;
		Dplus[62] = 18'b000000000_111100010;
		Dplus[63] = 18'b000000000_111100001;
		Dplus[64] = 18'b000000000_111100001;
		Dplus[65] = 18'b000000000_111100000;
		Dplus[66] = 18'b000000000_111100000;
		Dplus[67] = 18'b000000000_111011111;
		Dplus[68] = 18'b000000000_111011111;
		Dplus[69] = 18'b000000000_111011110;
		Dplus[70] = 18'b000000000_111011110;
		Dplus[71] = 18'b000000000_111011101;
		Dplus[72] = 18'b000000000_111011101;
		Dplus[73] = 18'b000000000_111011100;
		Dplus[74] = 18'b000000000_111011100;
		Dplus[75] = 18'b000000000_111011011;
		Dplus[76] = 18'b000000000_111011011;
		Dplus[77] = 18'b000000000_111011011;
		Dplus[78] = 18'b000000000_111011010;
		Dplus[79] = 18'b000000000_111011010;
		Dplus[80] = 18'b000000000_111011001;
		Dplus[81] = 18'b000000000_111011001;
		Dplus[82] = 18'b000000000_111011000;
		Dplus[83] = 18'b000000000_111011000;
		Dplus[84] = 18'b000000000_111010111;
		Dplus[85] = 18'b000000000_111010111;
		Dplus[86] = 18'b000000000_111010110;
		Dplus[87] = 18'b000000000_111010110;
		Dplus[88] = 18'b000000000_111010101;
		Dplus[89] = 18'b000000000_111010101;
		Dplus[90] = 18'b000000000_111010100;
		Dplus[91] = 18'b000000000_111010100;
		Dplus[92] = 18'b000000000_111010011;
		Dplus[93] = 18'b000000000_111010011;
		Dplus[94] = 18'b000000000_111010010;
		Dplus[95] = 18'b000000000_111010010;
		Dplus[96] = 18'b000000000_111010010;
		Dplus[97] = 18'b000000000_111010001;
		Dplus[98] = 18'b000000000_111010001;
		Dplus[99] = 18'b000000000_111010000;
		Dplus[100] = 18'b000000000_111010000;
		Dplus[101] = 18'b000000000_111001111;
		Dplus[102] = 18'b000000000_111001111;
		Dplus[103] = 18'b000000000_111001110;
		Dplus[104] = 18'b000000000_111001110;
		Dplus[105] = 18'b000000000_111001101;
		Dplus[106] = 18'b000000000_111001101;
		Dplus[107] = 18'b000000000_111001100;
		Dplus[108] = 18'b000000000_111001100;
		Dplus[109] = 18'b000000000_111001100;
		Dplus[110] = 18'b000000000_111001011;
		Dplus[111] = 18'b000000000_111001011;
		Dplus[112] = 18'b000000000_111001010;
		Dplus[113] = 18'b000000000_111001010;
		Dplus[114] = 18'b000000000_111001001;
		Dplus[115] = 18'b000000000_111001001;
		Dplus[116] = 18'b000000000_111001000;
		Dplus[117] = 18'b000000000_111001000;
		Dplus[118] = 18'b000000000_111000111;
		Dplus[119] = 18'b000000000_111000111;
		Dplus[120] = 18'b000000000_111000110;
		Dplus[121] = 18'b000000000_111000110;
		Dplus[122] = 18'b000000000_111000110;
		Dplus[123] = 18'b000000000_111000101;
		Dplus[124] = 18'b000000000_111000101;
		Dplus[125] = 18'b000000000_111000100;
		Dplus[126] = 18'b000000000_111000100;
		Dplus[127] = 18'b000000000_111000011;
		Dplus[128] = 18'b000000000_111000011;
		Dplus[129] = 18'b000000000_111000010;
		Dplus[130] = 18'b000000000_111000010;
		Dplus[131] = 18'b000000000_111000001;
		Dplus[132] = 18'b000000000_111000001;
		Dplus[133] = 18'b000000000_111000000;
		Dplus[134] = 18'b000000000_111000000;
		Dplus[135] = 18'b000000000_111000000;
		Dplus[136] = 18'b000000000_110111111;
		Dplus[137] = 18'b000000000_110111111;
		Dplus[138] = 18'b000000000_110111110;
		Dplus[139] = 18'b000000000_110111110;
		Dplus[140] = 18'b000000000_110111101;
		Dplus[141] = 18'b000000000_110111101;
		Dplus[142] = 18'b000000000_110111100;
		Dplus[143] = 18'b000000000_110111100;
		Dplus[144] = 18'b000000000_110111100;
		Dplus[145] = 18'b000000000_110111011;
		Dplus[146] = 18'b000000000_110111011;
		Dplus[147] = 18'b000000000_110111010;
		Dplus[148] = 18'b000000000_110111010;
		Dplus[149] = 18'b000000000_110111001;
		Dplus[150] = 18'b000000000_110111001;
		Dplus[151] = 18'b000000000_110111000;
		Dplus[152] = 18'b000000000_110111000;
		Dplus[153] = 18'b000000000_110110111;
		Dplus[154] = 18'b000000000_110110111;
		Dplus[155] = 18'b000000000_110110111;
		Dplus[156] = 18'b000000000_110110110;
		Dplus[157] = 18'b000000000_110110110;
		Dplus[158] = 18'b000000000_110110101;
		Dplus[159] = 18'b000000000_110110101;
		Dplus[160] = 18'b000000000_110110100;
		Dplus[161] = 18'b000000000_110110100;
		Dplus[162] = 18'b000000000_110110011;
		Dplus[163] = 18'b000000000_110110011;
		Dplus[164] = 18'b000000000_110110011;
		Dplus[165] = 18'b000000000_110110010;
		Dplus[166] = 18'b000000000_110110010;
		Dplus[167] = 18'b000000000_110110001;
		Dplus[168] = 18'b000000000_110110001;
		Dplus[169] = 18'b000000000_110110000;
		Dplus[170] = 18'b000000000_110110000;
		Dplus[171] = 18'b000000000_110101111;
		Dplus[172] = 18'b000000000_110101111;
		Dplus[173] = 18'b000000000_110101111;
		Dplus[174] = 18'b000000000_110101110;
		Dplus[175] = 18'b000000000_110101110;
		Dplus[176] = 18'b000000000_110101101;
		Dplus[177] = 18'b000000000_110101101;
		Dplus[178] = 18'b000000000_110101100;
		Dplus[179] = 18'b000000000_110101100;
		Dplus[180] = 18'b000000000_110101011;
		Dplus[181] = 18'b000000000_110101011;
		Dplus[182] = 18'b000000000_110101011;
		Dplus[183] = 18'b000000000_110101010;
		Dplus[184] = 18'b000000000_110101010;
		Dplus[185] = 18'b000000000_110101001;
		Dplus[186] = 18'b000000000_110101001;
		Dplus[187] = 18'b000000000_110101000;
		Dplus[188] = 18'b000000000_110101000;
		Dplus[189] = 18'b000000000_110101000;
		Dplus[190] = 18'b000000000_110100111;
		Dplus[191] = 18'b000000000_110100111;
		Dplus[192] = 18'b000000000_110100110;
		Dplus[193] = 18'b000000000_110100110;
		Dplus[194] = 18'b000000000_110100101;
		Dplus[195] = 18'b000000000_110100101;
		Dplus[196] = 18'b000000000_110100100;
		Dplus[197] = 18'b000000000_110100100;
		Dplus[198] = 18'b000000000_110100100;
		Dplus[199] = 18'b000000000_110100011;
		Dplus[200] = 18'b000000000_110100011;
		Dplus[201] = 18'b000000000_110100010;
		Dplus[202] = 18'b000000000_110100010;
		Dplus[203] = 18'b000000000_110100001;
		Dplus[204] = 18'b000000000_110100001;
		Dplus[205] = 18'b000000000_110100001;
		Dplus[206] = 18'b000000000_110100000;
		Dplus[207] = 18'b000000000_110100000;
		Dplus[208] = 18'b000000000_110011111;
		Dplus[209] = 18'b000000000_110011111;
		Dplus[210] = 18'b000000000_110011110;
		Dplus[211] = 18'b000000000_110011110;
		Dplus[212] = 18'b000000000_110011110;
		Dplus[213] = 18'b000000000_110011101;
		Dplus[214] = 18'b000000000_110011101;
		Dplus[215] = 18'b000000000_110011100;
		Dplus[216] = 18'b000000000_110011100;
		Dplus[217] = 18'b000000000_110011011;
		Dplus[218] = 18'b000000000_110011011;
		Dplus[219] = 18'b000000000_110011011;
		Dplus[220] = 18'b000000000_110011010;
		Dplus[221] = 18'b000000000_110011010;
		Dplus[222] = 18'b000000000_110011001;
		Dplus[223] = 18'b000000000_110011001;
		Dplus[224] = 18'b000000000_110011000;
		Dplus[225] = 18'b000000000_110011000;
		Dplus[226] = 18'b000000000_110011000;
		Dplus[227] = 18'b000000000_110010111;
		Dplus[228] = 18'b000000000_110010111;
		Dplus[229] = 18'b000000000_110010110;
		Dplus[230] = 18'b000000000_110010110;
		Dplus[231] = 18'b000000000_110010101;
		Dplus[232] = 18'b000000000_110010101;
		Dplus[233] = 18'b000000000_110010101;
		Dplus[234] = 18'b000000000_110010100;
		Dplus[235] = 18'b000000000_110010100;
		Dplus[236] = 18'b000000000_110010011;
		Dplus[237] = 18'b000000000_110010011;
		Dplus[238] = 18'b000000000_110010011;
		Dplus[239] = 18'b000000000_110010010;
		Dplus[240] = 18'b000000000_110010010;
		Dplus[241] = 18'b000000000_110010001;
		Dplus[242] = 18'b000000000_110010001;
		Dplus[243] = 18'b000000000_110010000;
		Dplus[244] = 18'b000000000_110010000;
		Dplus[245] = 18'b000000000_110010000;
		Dplus[246] = 18'b000000000_110001111;
		Dplus[247] = 18'b000000000_110001111;
		Dplus[248] = 18'b000000000_110001110;
		Dplus[249] = 18'b000000000_110001110;
		Dplus[250] = 18'b000000000_110001110;
		Dplus[251] = 18'b000000000_110001101;
		Dplus[252] = 18'b000000000_110001101;
		Dplus[253] = 18'b000000000_110001100;
		Dplus[254] = 18'b000000000_110001100;
		Dplus[255] = 18'b000000000_110001011;
		Dplus[256] = 18'b000000000_110001011;
		Dplus[257] = 18'b000000000_110001011;
		Dplus[258] = 18'b000000000_110001010;
		Dplus[259] = 18'b000000000_110001010;
		Dplus[260] = 18'b000000000_110001001;
		Dplus[261] = 18'b000000000_110001001;
		Dplus[262] = 18'b000000000_110001001;
		Dplus[263] = 18'b000000000_110001000;
		Dplus[264] = 18'b000000000_110001000;
		Dplus[265] = 18'b000000000_110000111;
		Dplus[266] = 18'b000000000_110000111;
		Dplus[267] = 18'b000000000_110000110;
		Dplus[268] = 18'b000000000_110000110;
		Dplus[269] = 18'b000000000_110000110;
		Dplus[270] = 18'b000000000_110000101;
		Dplus[271] = 18'b000000000_110000101;
		Dplus[272] = 18'b000000000_110000100;
		Dplus[273] = 18'b000000000_110000100;
		Dplus[274] = 18'b000000000_110000100;
		Dplus[275] = 18'b000000000_110000011;
		Dplus[276] = 18'b000000000_110000011;
		Dplus[277] = 18'b000000000_110000010;
		Dplus[278] = 18'b000000000_110000010;
		Dplus[279] = 18'b000000000_110000010;
		Dplus[280] = 18'b000000000_110000001;
		Dplus[281] = 18'b000000000_110000001;
		Dplus[282] = 18'b000000000_110000000;
		Dplus[283] = 18'b000000000_110000000;
		Dplus[284] = 18'b000000000_110000000;
		Dplus[285] = 18'b000000000_101111111;
		Dplus[286] = 18'b000000000_101111111;
		Dplus[287] = 18'b000000000_101111110;
		Dplus[288] = 18'b000000000_101111110;
		Dplus[289] = 18'b000000000_101111110;
		Dplus[290] = 18'b000000000_101111101;
		Dplus[291] = 18'b000000000_101111101;
		Dplus[292] = 18'b000000000_101111100;
		Dplus[293] = 18'b000000000_101111100;
		Dplus[294] = 18'b000000000_101111100;
		Dplus[295] = 18'b000000000_101111011;
		Dplus[296] = 18'b000000000_101111011;
		Dplus[297] = 18'b000000000_101111010;
		Dplus[298] = 18'b000000000_101111010;
		Dplus[299] = 18'b000000000_101111010;
		Dplus[300] = 18'b000000000_101111001;
		Dplus[301] = 18'b000000000_101111001;
		Dplus[302] = 18'b000000000_101111000;
		Dplus[303] = 18'b000000000_101111000;
		Dplus[304] = 18'b000000000_101111000;
		Dplus[305] = 18'b000000000_101110111;
		Dplus[306] = 18'b000000000_101110111;
		Dplus[307] = 18'b000000000_101110110;
		Dplus[308] = 18'b000000000_101110110;
		Dplus[309] = 18'b000000000_101110110;
		Dplus[310] = 18'b000000000_101110101;
		Dplus[311] = 18'b000000000_101110101;
		Dplus[312] = 18'b000000000_101110100;
		Dplus[313] = 18'b000000000_101110100;
		Dplus[314] = 18'b000000000_101110100;
		Dplus[315] = 18'b000000000_101110011;
		Dplus[316] = 18'b000000000_101110011;
		Dplus[317] = 18'b000000000_101110010;
		Dplus[318] = 18'b000000000_101110010;
		Dplus[319] = 18'b000000000_101110010;
		Dplus[320] = 18'b000000000_101110001;
		Dplus[321] = 18'b000000000_101110001;
		Dplus[322] = 18'b000000000_101110000;
		Dplus[323] = 18'b000000000_101110000;
		Dplus[324] = 18'b000000000_101110000;
		Dplus[325] = 18'b000000000_101101111;
		Dplus[326] = 18'b000000000_101101111;
		Dplus[327] = 18'b000000000_101101110;
		Dplus[328] = 18'b000000000_101101110;
		Dplus[329] = 18'b000000000_101101110;
		Dplus[330] = 18'b000000000_101101101;
		Dplus[331] = 18'b000000000_101101101;
		Dplus[332] = 18'b000000000_101101100;
		Dplus[333] = 18'b000000000_101101100;
		Dplus[334] = 18'b000000000_101101100;
		Dplus[335] = 18'b000000000_101101011;
		Dplus[336] = 18'b000000000_101101011;
		Dplus[337] = 18'b000000000_101101011;
		Dplus[338] = 18'b000000000_101101010;
		Dplus[339] = 18'b000000000_101101010;
		Dplus[340] = 18'b000000000_101101001;
		Dplus[341] = 18'b000000000_101101001;
		Dplus[342] = 18'b000000000_101101001;
		Dplus[343] = 18'b000000000_101101000;
		Dplus[344] = 18'b000000000_101101000;
		Dplus[345] = 18'b000000000_101100111;
		Dplus[346] = 18'b000000000_101100111;
		Dplus[347] = 18'b000000000_101100111;
		Dplus[348] = 18'b000000000_101100110;
		Dplus[349] = 18'b000000000_101100110;
		Dplus[350] = 18'b000000000_101100110;
		Dplus[351] = 18'b000000000_101100101;
		Dplus[352] = 18'b000000000_101100101;
		Dplus[353] = 18'b000000000_101100100;
		Dplus[354] = 18'b000000000_101100100;
		Dplus[355] = 18'b000000000_101100100;
		Dplus[356] = 18'b000000000_101100011;
		Dplus[357] = 18'b000000000_101100011;
		Dplus[358] = 18'b000000000_101100010;
		Dplus[359] = 18'b000000000_101100010;
		Dplus[360] = 18'b000000000_101100010;
		Dplus[361] = 18'b000000000_101100001;
		Dplus[362] = 18'b000000000_101100001;
		Dplus[363] = 18'b000000000_101100001;
		Dplus[364] = 18'b000000000_101100000;
		Dplus[365] = 18'b000000000_101100000;
		Dplus[366] = 18'b000000000_101011111;
		Dplus[367] = 18'b000000000_101011111;
		Dplus[368] = 18'b000000000_101011111;
		Dplus[369] = 18'b000000000_101011110;
		Dplus[370] = 18'b000000000_101011110;
		Dplus[371] = 18'b000000000_101011110;
		Dplus[372] = 18'b000000000_101011101;
		Dplus[373] = 18'b000000000_101011101;
		Dplus[374] = 18'b000000000_101011100;
		Dplus[375] = 18'b000000000_101011100;
		Dplus[376] = 18'b000000000_101011100;
		Dplus[377] = 18'b000000000_101011011;
		Dplus[378] = 18'b000000000_101011011;
		Dplus[379] = 18'b000000000_101011011;
		Dplus[380] = 18'b000000000_101011010;
		Dplus[381] = 18'b000000000_101011010;
		Dplus[382] = 18'b000000000_101011001;
		Dplus[383] = 18'b000000000_101011001;
		Dplus[384] = 18'b000000000_101011001;
		Dplus[385] = 18'b000000000_101011000;
		Dplus[386] = 18'b000000000_101011000;
		Dplus[387] = 18'b000000000_101011000;
		Dplus[388] = 18'b000000000_101010111;
		Dplus[389] = 18'b000000000_101010111;
		Dplus[390] = 18'b000000000_101010110;
		Dplus[391] = 18'b000000000_101010110;
		Dplus[392] = 18'b000000000_101010110;
		Dplus[393] = 18'b000000000_101010101;
		Dplus[394] = 18'b000000000_101010101;
		Dplus[395] = 18'b000000000_101010101;
		Dplus[396] = 18'b000000000_101010100;
		Dplus[397] = 18'b000000000_101010100;
		Dplus[398] = 18'b000000000_101010011;
		Dplus[399] = 18'b000000000_101010011;
		Dplus[400] = 18'b000000000_101010011;
		Dplus[401] = 18'b000000000_101010010;
		Dplus[402] = 18'b000000000_101010010;
		Dplus[403] = 18'b000000000_101010010;
		Dplus[404] = 18'b000000000_101010001;
		Dplus[405] = 18'b000000000_101010001;
		Dplus[406] = 18'b000000000_101010001;
		Dplus[407] = 18'b000000000_101010000;
		Dplus[408] = 18'b000000000_101010000;
		Dplus[409] = 18'b000000000_101001111;
		Dplus[410] = 18'b000000000_101001111;
		Dplus[411] = 18'b000000000_101001111;
		Dplus[412] = 18'b000000000_101001110;
		Dplus[413] = 18'b000000000_101001110;
		Dplus[414] = 18'b000000000_101001110;
		Dplus[415] = 18'b000000000_101001101;
		Dplus[416] = 18'b000000000_101001101;
		Dplus[417] = 18'b000000000_101001101;
		Dplus[418] = 18'b000000000_101001100;
		Dplus[419] = 18'b000000000_101001100;
		Dplus[420] = 18'b000000000_101001011;
		Dplus[421] = 18'b000000000_101001011;
		Dplus[422] = 18'b000000000_101001011;
		Dplus[423] = 18'b000000000_101001010;
		Dplus[424] = 18'b000000000_101001010;
		Dplus[425] = 18'b000000000_101001010;
		Dplus[426] = 18'b000000000_101001001;
		Dplus[427] = 18'b000000000_101001001;
		Dplus[428] = 18'b000000000_101001001;
		Dplus[429] = 18'b000000000_101001000;
		Dplus[430] = 18'b000000000_101001000;
		Dplus[431] = 18'b000000000_101000111;
		Dplus[432] = 18'b000000000_101000111;
		Dplus[433] = 18'b000000000_101000111;
		Dplus[434] = 18'b000000000_101000110;
		Dplus[435] = 18'b000000000_101000110;
		Dplus[436] = 18'b000000000_101000110;
		Dplus[437] = 18'b000000000_101000101;
		Dplus[438] = 18'b000000000_101000101;
		Dplus[439] = 18'b000000000_101000101;
		Dplus[440] = 18'b000000000_101000100;
		Dplus[441] = 18'b000000000_101000100;
		Dplus[442] = 18'b000000000_101000100;
		Dplus[443] = 18'b000000000_101000011;
		Dplus[444] = 18'b000000000_101000011;
		Dplus[445] = 18'b000000000_101000011;
		Dplus[446] = 18'b000000000_101000010;
		Dplus[447] = 18'b000000000_101000010;
		Dplus[448] = 18'b000000000_101000001;
		Dplus[449] = 18'b000000000_101000001;
		Dplus[450] = 18'b000000000_101000001;
		Dplus[451] = 18'b000000000_101000000;
		Dplus[452] = 18'b000000000_101000000;
		Dplus[453] = 18'b000000000_101000000;
		Dplus[454] = 18'b000000000_100111111;
		Dplus[455] = 18'b000000000_100111111;
		Dplus[456] = 18'b000000000_100111111;
		Dplus[457] = 18'b000000000_100111110;
		Dplus[458] = 18'b000000000_100111110;
		Dplus[459] = 18'b000000000_100111110;
		Dplus[460] = 18'b000000000_100111101;
		Dplus[461] = 18'b000000000_100111101;
		Dplus[462] = 18'b000000000_100111101;
		Dplus[463] = 18'b000000000_100111100;
		Dplus[464] = 18'b000000000_100111100;
		Dplus[465] = 18'b000000000_100111100;
		Dplus[466] = 18'b000000000_100111011;
		Dplus[467] = 18'b000000000_100111011;
		Dplus[468] = 18'b000000000_100111010;
		Dplus[469] = 18'b000000000_100111010;
		Dplus[470] = 18'b000000000_100111010;
		Dplus[471] = 18'b000000000_100111001;
		Dplus[472] = 18'b000000000_100111001;
		Dplus[473] = 18'b000000000_100111001;
		Dplus[474] = 18'b000000000_100111000;
		Dplus[475] = 18'b000000000_100111000;
		Dplus[476] = 18'b000000000_100111000;
		Dplus[477] = 18'b000000000_100110111;
		Dplus[478] = 18'b000000000_100110111;
		Dplus[479] = 18'b000000000_100110111;
		Dplus[480] = 18'b000000000_100110110;
		Dplus[481] = 18'b000000000_100110110;
		Dplus[482] = 18'b000000000_100110110;
		Dplus[483] = 18'b000000000_100110101;
		Dplus[484] = 18'b000000000_100110101;
		Dplus[485] = 18'b000000000_100110101;
		Dplus[486] = 18'b000000000_100110100;
		Dplus[487] = 18'b000000000_100110100;
		Dplus[488] = 18'b000000000_100110100;
		Dplus[489] = 18'b000000000_100110011;
		Dplus[490] = 18'b000000000_100110011;
		Dplus[491] = 18'b000000000_100110011;
		Dplus[492] = 18'b000000000_100110010;
		Dplus[493] = 18'b000000000_100110010;
		Dplus[494] = 18'b000000000_100110010;
		Dplus[495] = 18'b000000000_100110001;
		Dplus[496] = 18'b000000000_100110001;
		Dplus[497] = 18'b000000000_100110001;
		Dplus[498] = 18'b000000000_100110000;
		Dplus[499] = 18'b000000000_100110000;
		Dplus[500] = 18'b000000000_100110000;
		Dplus[501] = 18'b000000000_100101111;
		Dplus[502] = 18'b000000000_100101111;
		Dplus[503] = 18'b000000000_100101111;
		Dplus[504] = 18'b000000000_100101110;
		Dplus[505] = 18'b000000000_100101110;
		Dplus[506] = 18'b000000000_100101110;
		Dplus[507] = 18'b000000000_100101101;
		Dplus[508] = 18'b000000000_100101101;
		Dplus[509] = 18'b000000000_100101101;
		Dplus[510] = 18'b000000000_100101100;
		Dplus[511] = 18'b000000000_100101100;
		Dplus[512] = 18'b000000000_100101100;
		Dplus[513] = 18'b000000000_100101011;
		Dplus[514] = 18'b000000000_100101011;
		Dplus[515] = 18'b000000000_100101011;
		Dplus[516] = 18'b000000000_100101010;
		Dplus[517] = 18'b000000000_100101010;
		Dplus[518] = 18'b000000000_100101010;
		Dplus[519] = 18'b000000000_100101001;
		Dplus[520] = 18'b000000000_100101001;
		Dplus[521] = 18'b000000000_100101001;
		Dplus[522] = 18'b000000000_100101000;
		Dplus[523] = 18'b000000000_100101000;
		Dplus[524] = 18'b000000000_100101000;
		Dplus[525] = 18'b000000000_100100111;
		Dplus[526] = 18'b000000000_100100111;
		Dplus[527] = 18'b000000000_100100111;
		Dplus[528] = 18'b000000000_100100110;
		Dplus[529] = 18'b000000000_100100110;
		Dplus[530] = 18'b000000000_100100110;
		Dplus[531] = 18'b000000000_100100101;
		Dplus[532] = 18'b000000000_100100101;
		Dplus[533] = 18'b000000000_100100101;
		Dplus[534] = 18'b000000000_100100100;
		Dplus[535] = 18'b000000000_100100100;
		Dplus[536] = 18'b000000000_100100100;
		Dplus[537] = 18'b000000000_100100011;
		Dplus[538] = 18'b000000000_100100011;
		Dplus[539] = 18'b000000000_100100011;
		Dplus[540] = 18'b000000000_100100010;
		Dplus[541] = 18'b000000000_100100010;
		Dplus[542] = 18'b000000000_100100010;
		Dplus[543] = 18'b000000000_100100001;
		Dplus[544] = 18'b000000000_100100001;
		Dplus[545] = 18'b000000000_100100001;
		Dplus[546] = 18'b000000000_100100000;
		Dplus[547] = 18'b000000000_100100000;
		Dplus[548] = 18'b000000000_100100000;
		Dplus[549] = 18'b000000000_100011111;
		Dplus[550] = 18'b000000000_100011111;
		Dplus[551] = 18'b000000000_100011111;
		Dplus[552] = 18'b000000000_100011110;
		Dplus[553] = 18'b000000000_100011110;
		Dplus[554] = 18'b000000000_100011110;
		Dplus[555] = 18'b000000000_100011101;
		Dplus[556] = 18'b000000000_100011101;
		Dplus[557] = 18'b000000000_100011101;
		Dplus[558] = 18'b000000000_100011100;
		Dplus[559] = 18'b000000000_100011100;
		Dplus[560] = 18'b000000000_100011100;
		Dplus[561] = 18'b000000000_100011100;
		Dplus[562] = 18'b000000000_100011011;
		Dplus[563] = 18'b000000000_100011011;
		Dplus[564] = 18'b000000000_100011011;
		Dplus[565] = 18'b000000000_100011010;
		Dplus[566] = 18'b000000000_100011010;
		Dplus[567] = 18'b000000000_100011010;
		Dplus[568] = 18'b000000000_100011001;
		Dplus[569] = 18'b000000000_100011001;
		Dplus[570] = 18'b000000000_100011001;
		Dplus[571] = 18'b000000000_100011000;
		Dplus[572] = 18'b000000000_100011000;
		Dplus[573] = 18'b000000000_100011000;
		Dplus[574] = 18'b000000000_100010111;
		Dplus[575] = 18'b000000000_100010111;
		Dplus[576] = 18'b000000000_100010111;
		Dplus[577] = 18'b000000000_100010110;
		Dplus[578] = 18'b000000000_100010110;
		Dplus[579] = 18'b000000000_100010110;
		Dplus[580] = 18'b000000000_100010110;
		Dplus[581] = 18'b000000000_100010101;
		Dplus[582] = 18'b000000000_100010101;
		Dplus[583] = 18'b000000000_100010101;
		Dplus[584] = 18'b000000000_100010100;
		Dplus[585] = 18'b000000000_100010100;
		Dplus[586] = 18'b000000000_100010100;
		Dplus[587] = 18'b000000000_100010011;
		Dplus[588] = 18'b000000000_100010011;
		Dplus[589] = 18'b000000000_100010011;
		Dplus[590] = 18'b000000000_100010010;
		Dplus[591] = 18'b000000000_100010010;
		Dplus[592] = 18'b000000000_100010010;
		Dplus[593] = 18'b000000000_100010001;
		Dplus[594] = 18'b000000000_100010001;
		Dplus[595] = 18'b000000000_100010001;
		Dplus[596] = 18'b000000000_100010001;
		Dplus[597] = 18'b000000000_100010000;
		Dplus[598] = 18'b000000000_100010000;
		Dplus[599] = 18'b000000000_100010000;
		Dplus[600] = 18'b000000000_100001111;
		Dplus[601] = 18'b000000000_100001111;
		Dplus[602] = 18'b000000000_100001111;
		Dplus[603] = 18'b000000000_100001110;
		Dplus[604] = 18'b000000000_100001110;
		Dplus[605] = 18'b000000000_100001110;
		Dplus[606] = 18'b000000000_100001101;
		Dplus[607] = 18'b000000000_100001101;
		Dplus[608] = 18'b000000000_100001101;
		Dplus[609] = 18'b000000000_100001101;
		Dplus[610] = 18'b000000000_100001100;
		Dplus[611] = 18'b000000000_100001100;
		Dplus[612] = 18'b000000000_100001100;
		Dplus[613] = 18'b000000000_100001011;
		Dplus[614] = 18'b000000000_100001011;
		Dplus[615] = 18'b000000000_100001011;
		Dplus[616] = 18'b000000000_100001010;
		Dplus[617] = 18'b000000000_100001010;
		Dplus[618] = 18'b000000000_100001010;
		Dplus[619] = 18'b000000000_100001010;
		Dplus[620] = 18'b000000000_100001001;
		Dplus[621] = 18'b000000000_100001001;
		Dplus[622] = 18'b000000000_100001001;
		Dplus[623] = 18'b000000000_100001000;
		Dplus[624] = 18'b000000000_100001000;
		Dplus[625] = 18'b000000000_100001000;
		Dplus[626] = 18'b000000000_100000111;
		Dplus[627] = 18'b000000000_100000111;
		Dplus[628] = 18'b000000000_100000111;
		Dplus[629] = 18'b000000000_100000111;
		Dplus[630] = 18'b000000000_100000110;
		Dplus[631] = 18'b000000000_100000110;
		Dplus[632] = 18'b000000000_100000110;
		Dplus[633] = 18'b000000000_100000101;
		Dplus[634] = 18'b000000000_100000101;
		Dplus[635] = 18'b000000000_100000101;
		Dplus[636] = 18'b000000000_100000100;
		Dplus[637] = 18'b000000000_100000100;
		Dplus[638] = 18'b000000000_100000100;
		Dplus[639] = 18'b000000000_100000100;
		Dplus[640] = 18'b000000000_100000011;
		Dplus[641] = 18'b000000000_100000011;
		Dplus[642] = 18'b000000000_100000011;
		Dplus[643] = 18'b000000000_100000010;
		Dplus[644] = 18'b000000000_100000010;
		Dplus[645] = 18'b000000000_100000010;
		Dplus[646] = 18'b000000000_100000001;
		Dplus[647] = 18'b000000000_100000001;
		Dplus[648] = 18'b000000000_100000001;
		Dplus[649] = 18'b000000000_100000001;
		Dplus[650] = 18'b000000000_100000000;
		Dplus[651] = 18'b000000000_100000000;
		Dplus[652] = 18'b000000000_100000000;
		Dplus[653] = 18'b000000000_011111111;
		Dplus[654] = 18'b000000000_011111111;
		Dplus[655] = 18'b000000000_011111111;
		Dplus[656] = 18'b000000000_011111111;
		Dplus[657] = 18'b000000000_011111110;
		Dplus[658] = 18'b000000000_011111110;
		Dplus[659] = 18'b000000000_011111110;
		Dplus[660] = 18'b000000000_011111101;
		Dplus[661] = 18'b000000000_011111101;
		Dplus[662] = 18'b000000000_011111101;
		Dplus[663] = 18'b000000000_011111101;
		Dplus[664] = 18'b000000000_011111100;
		Dplus[665] = 18'b000000000_011111100;
		Dplus[666] = 18'b000000000_011111100;
		Dplus[667] = 18'b000000000_011111011;
		Dplus[668] = 18'b000000000_011111011;
		Dplus[669] = 18'b000000000_011111011;
		Dplus[670] = 18'b000000000_011111010;
		Dplus[671] = 18'b000000000_011111010;
		Dplus[672] = 18'b000000000_011111010;
		Dplus[673] = 18'b000000000_011111010;
		Dplus[674] = 18'b000000000_011111001;
		Dplus[675] = 18'b000000000_011111001;
		Dplus[676] = 18'b000000000_011111001;
		Dplus[677] = 18'b000000000_011111000;
		Dplus[678] = 18'b000000000_011111000;
		Dplus[679] = 18'b000000000_011111000;
		Dplus[680] = 18'b000000000_011111000;
		Dplus[681] = 18'b000000000_011110111;
		Dplus[682] = 18'b000000000_011110111;
		Dplus[683] = 18'b000000000_011110111;
		Dplus[684] = 18'b000000000_011110110;
		Dplus[685] = 18'b000000000_011110110;
		Dplus[686] = 18'b000000000_011110110;
		Dplus[687] = 18'b000000000_011110110;
		Dplus[688] = 18'b000000000_011110101;
		Dplus[689] = 18'b000000000_011110101;
		Dplus[690] = 18'b000000000_011110101;
		Dplus[691] = 18'b000000000_011110101;
		Dplus[692] = 18'b000000000_011110100;
		Dplus[693] = 18'b000000000_011110100;
		Dplus[694] = 18'b000000000_011110100;
		Dplus[695] = 18'b000000000_011110011;
		Dplus[696] = 18'b000000000_011110011;
		Dplus[697] = 18'b000000000_011110011;
		Dplus[698] = 18'b000000000_011110011;
		Dplus[699] = 18'b000000000_011110010;
		Dplus[700] = 18'b000000000_011110010;
		Dplus[701] = 18'b000000000_011110010;
		Dplus[702] = 18'b000000000_011110001;
		Dplus[703] = 18'b000000000_011110001;
		Dplus[704] = 18'b000000000_011110001;
		Dplus[705] = 18'b000000000_011110001;
		Dplus[706] = 18'b000000000_011110000;
		Dplus[707] = 18'b000000000_011110000;
		Dplus[708] = 18'b000000000_011110000;
		Dplus[709] = 18'b000000000_011101111;
		Dplus[710] = 18'b000000000_011101111;
		Dplus[711] = 18'b000000000_011101111;
		Dplus[712] = 18'b000000000_011101111;
		Dplus[713] = 18'b000000000_011101110;
		Dplus[714] = 18'b000000000_011101110;
		Dplus[715] = 18'b000000000_011101110;
		Dplus[716] = 18'b000000000_011101110;
		Dplus[717] = 18'b000000000_011101101;
		Dplus[718] = 18'b000000000_011101101;
		Dplus[719] = 18'b000000000_011101101;
		Dplus[720] = 18'b000000000_011101100;
		Dplus[721] = 18'b000000000_011101100;
		Dplus[722] = 18'b000000000_011101100;
		Dplus[723] = 18'b000000000_011101100;
		Dplus[724] = 18'b000000000_011101011;
		Dplus[725] = 18'b000000000_011101011;
		Dplus[726] = 18'b000000000_011101011;
		Dplus[727] = 18'b000000000_011101011;
		Dplus[728] = 18'b000000000_011101010;
		Dplus[729] = 18'b000000000_011101010;
		Dplus[730] = 18'b000000000_011101010;
		Dplus[731] = 18'b000000000_011101001;
		Dplus[732] = 18'b000000000_011101001;
		Dplus[733] = 18'b000000000_011101001;
		Dplus[734] = 18'b000000000_011101001;
		Dplus[735] = 18'b000000000_011101000;
		Dplus[736] = 18'b000000000_011101000;
		Dplus[737] = 18'b000000000_011101000;
		Dplus[738] = 18'b000000000_011101000;
		Dplus[739] = 18'b000000000_011100111;
		Dplus[740] = 18'b000000000_011100111;
		Dplus[741] = 18'b000000000_011100111;
		Dplus[742] = 18'b000000000_011100110;
		Dplus[743] = 18'b000000000_011100110;
		Dplus[744] = 18'b000000000_011100110;
		Dplus[745] = 18'b000000000_011100110;
		Dplus[746] = 18'b000000000_011100101;
		Dplus[747] = 18'b000000000_011100101;
		Dplus[748] = 18'b000000000_011100101;
		Dplus[749] = 18'b000000000_011100101;
		Dplus[750] = 18'b000000000_011100100;
		Dplus[751] = 18'b000000000_011100100;
		Dplus[752] = 18'b000000000_011100100;
		Dplus[753] = 18'b000000000_011100100;
		Dplus[754] = 18'b000000000_011100011;
		Dplus[755] = 18'b000000000_011100011;
		Dplus[756] = 18'b000000000_011100011;
		Dplus[757] = 18'b000000000_011100011;
		Dplus[758] = 18'b000000000_011100010;
		Dplus[759] = 18'b000000000_011100010;
		Dplus[760] = 18'b000000000_011100010;
		Dplus[761] = 18'b000000000_011100001;
		Dplus[762] = 18'b000000000_011100001;
		Dplus[763] = 18'b000000000_011100001;
		Dplus[764] = 18'b000000000_011100001;
		Dplus[765] = 18'b000000000_011100000;
		Dplus[766] = 18'b000000000_011100000;
		Dplus[767] = 18'b000000000_011100000;
		Dplus[768] = 18'b000000000_011100000;
		Dplus[769] = 18'b000000000_011011111;
		Dplus[770] = 18'b000000000_011011111;
		Dplus[771] = 18'b000000000_011011111;
		Dplus[772] = 18'b000000000_011011111;
		Dplus[773] = 18'b000000000_011011110;
		Dplus[774] = 18'b000000000_011011110;
		Dplus[775] = 18'b000000000_011011110;
		Dplus[776] = 18'b000000000_011011110;
		Dplus[777] = 18'b000000000_011011101;
		Dplus[778] = 18'b000000000_011011101;
		Dplus[779] = 18'b000000000_011011101;
		Dplus[780] = 18'b000000000_011011101;
		Dplus[781] = 18'b000000000_011011100;
		Dplus[782] = 18'b000000000_011011100;
		Dplus[783] = 18'b000000000_011011100;
		Dplus[784] = 18'b000000000_011011011;
		Dplus[785] = 18'b000000000_011011011;
		Dplus[786] = 18'b000000000_011011011;
		Dplus[787] = 18'b000000000_011011011;
		Dplus[788] = 18'b000000000_011011010;
		Dplus[789] = 18'b000000000_011011010;
		Dplus[790] = 18'b000000000_011011010;
		Dplus[791] = 18'b000000000_011011010;
		Dplus[792] = 18'b000000000_011011001;
		Dplus[793] = 18'b000000000_011011001;
		Dplus[794] = 18'b000000000_011011001;
		Dplus[795] = 18'b000000000_011011001;
		Dplus[796] = 18'b000000000_011011000;
		Dplus[797] = 18'b000000000_011011000;
		Dplus[798] = 18'b000000000_011011000;
		Dplus[799] = 18'b000000000_011011000;
		Dplus[800] = 18'b000000000_011010111;
		Dplus[801] = 18'b000000000_011010111;
		Dplus[802] = 18'b000000000_011010111;
		Dplus[803] = 18'b000000000_011010111;
		Dplus[804] = 18'b000000000_011010110;
		Dplus[805] = 18'b000000000_011010110;
		Dplus[806] = 18'b000000000_011010110;
		Dplus[807] = 18'b000000000_011010110;
		Dplus[808] = 18'b000000000_011010101;
		Dplus[809] = 18'b000000000_011010101;
		Dplus[810] = 18'b000000000_011010101;
		Dplus[811] = 18'b000000000_011010101;
		Dplus[812] = 18'b000000000_011010100;
		Dplus[813] = 18'b000000000_011010100;
		Dplus[814] = 18'b000000000_011010100;
		Dplus[815] = 18'b000000000_011010100;
		Dplus[816] = 18'b000000000_011010011;
		Dplus[817] = 18'b000000000_011010011;
		Dplus[818] = 18'b000000000_011010011;
		Dplus[819] = 18'b000000000_011010011;
		Dplus[820] = 18'b000000000_011010010;
		Dplus[821] = 18'b000000000_011010010;
		Dplus[822] = 18'b000000000_011010010;
		Dplus[823] = 18'b000000000_011010010;
		Dplus[824] = 18'b000000000_011010001;
		Dplus[825] = 18'b000000000_011010001;
		Dplus[826] = 18'b000000000_011010001;
		Dplus[827] = 18'b000000000_011010001;
		Dplus[828] = 18'b000000000_011010000;
		Dplus[829] = 18'b000000000_011010000;
		Dplus[830] = 18'b000000000_011010000;
		Dplus[831] = 18'b000000000_011010000;
		Dplus[832] = 18'b000000000_011001111;
		Dplus[833] = 18'b000000000_011001111;
		Dplus[834] = 18'b000000000_011001111;
		Dplus[835] = 18'b000000000_011001111;
		Dplus[836] = 18'b000000000_011001110;
		Dplus[837] = 18'b000000000_011001110;
		Dplus[838] = 18'b000000000_011001110;
		Dplus[839] = 18'b000000000_011001110;
		Dplus[840] = 18'b000000000_011001101;
		Dplus[841] = 18'b000000000_011001101;
		Dplus[842] = 18'b000000000_011001101;
		Dplus[843] = 18'b000000000_011001101;
		Dplus[844] = 18'b000000000_011001101;
		Dplus[845] = 18'b000000000_011001100;
		Dplus[846] = 18'b000000000_011001100;
		Dplus[847] = 18'b000000000_011001100;
		Dplus[848] = 18'b000000000_011001100;
		Dplus[849] = 18'b000000000_011001011;
		Dplus[850] = 18'b000000000_011001011;
		Dplus[851] = 18'b000000000_011001011;
		Dplus[852] = 18'b000000000_011001011;
		Dplus[853] = 18'b000000000_011001010;
		Dplus[854] = 18'b000000000_011001010;
		Dplus[855] = 18'b000000000_011001010;
		Dplus[856] = 18'b000000000_011001010;
		Dplus[857] = 18'b000000000_011001001;
		Dplus[858] = 18'b000000000_011001001;
		Dplus[859] = 18'b000000000_011001001;
		Dplus[860] = 18'b000000000_011001001;
		Dplus[861] = 18'b000000000_011001000;
		Dplus[862] = 18'b000000000_011001000;
		Dplus[863] = 18'b000000000_011001000;
		Dplus[864] = 18'b000000000_011001000;
		Dplus[865] = 18'b000000000_011000111;
		Dplus[866] = 18'b000000000_011000111;
		Dplus[867] = 18'b000000000_011000111;
		Dplus[868] = 18'b000000000_011000111;
		Dplus[869] = 18'b000000000_011000111;
		Dplus[870] = 18'b000000000_011000110;
		Dplus[871] = 18'b000000000_011000110;
		Dplus[872] = 18'b000000000_011000110;
		Dplus[873] = 18'b000000000_011000110;
		Dplus[874] = 18'b000000000_011000101;
		Dplus[875] = 18'b000000000_011000101;
		Dplus[876] = 18'b000000000_011000101;
		Dplus[877] = 18'b000000000_011000101;
		Dplus[878] = 18'b000000000_011000100;
		Dplus[879] = 18'b000000000_011000100;
		Dplus[880] = 18'b000000000_011000100;
		Dplus[881] = 18'b000000000_011000100;
		Dplus[882] = 18'b000000000_011000011;
		Dplus[883] = 18'b000000000_011000011;
		Dplus[884] = 18'b000000000_011000011;
		Dplus[885] = 18'b000000000_011000011;
		Dplus[886] = 18'b000000000_011000011;
		Dplus[887] = 18'b000000000_011000010;
		Dplus[888] = 18'b000000000_011000010;
		Dplus[889] = 18'b000000000_011000010;
		Dplus[890] = 18'b000000000_011000010;
		Dplus[891] = 18'b000000000_011000001;
		Dplus[892] = 18'b000000000_011000001;
		Dplus[893] = 18'b000000000_011000001;
		Dplus[894] = 18'b000000000_011000001;
		Dplus[895] = 18'b000000000_011000000;
		Dplus[896] = 18'b000000000_011000000;
		Dplus[897] = 18'b000000000_011000000;
		Dplus[898] = 18'b000000000_011000000;
		Dplus[899] = 18'b000000000_011000000;
		Dplus[900] = 18'b000000000_010111111;
		Dplus[901] = 18'b000000000_010111111;
		Dplus[902] = 18'b000000000_010111111;
		Dplus[903] = 18'b000000000_010111111;
		Dplus[904] = 18'b000000000_010111110;
		Dplus[905] = 18'b000000000_010111110;
		Dplus[906] = 18'b000000000_010111110;
		Dplus[907] = 18'b000000000_010111110;
		Dplus[908] = 18'b000000000_010111110;
		Dplus[909] = 18'b000000000_010111101;
		Dplus[910] = 18'b000000000_010111101;
		Dplus[911] = 18'b000000000_010111101;
		Dplus[912] = 18'b000000000_010111101;
		Dplus[913] = 18'b000000000_010111100;
		Dplus[914] = 18'b000000000_010111100;
		Dplus[915] = 18'b000000000_010111100;
		Dplus[916] = 18'b000000000_010111100;
		Dplus[917] = 18'b000000000_010111100;
		Dplus[918] = 18'b000000000_010111011;
		Dplus[919] = 18'b000000000_010111011;
		Dplus[920] = 18'b000000000_010111011;
		Dplus[921] = 18'b000000000_010111011;
		Dplus[922] = 18'b000000000_010111010;
		Dplus[923] = 18'b000000000_010111010;
		Dplus[924] = 18'b000000000_010111010;
		Dplus[925] = 18'b000000000_010111010;
		Dplus[926] = 18'b000000000_010111001;
		Dplus[927] = 18'b000000000_010111001;
		Dplus[928] = 18'b000000000_010111001;
		Dplus[929] = 18'b000000000_010111001;
		Dplus[930] = 18'b000000000_010111001;
		Dplus[931] = 18'b000000000_010111000;
		Dplus[932] = 18'b000000000_010111000;
		Dplus[933] = 18'b000000000_010111000;
		Dplus[934] = 18'b000000000_010111000;
		Dplus[935] = 18'b000000000_010111000;
		Dplus[936] = 18'b000000000_010110111;
		Dplus[937] = 18'b000000000_010110111;
		Dplus[938] = 18'b000000000_010110111;
		Dplus[939] = 18'b000000000_010110111;
		Dplus[940] = 18'b000000000_010110110;
		Dplus[941] = 18'b000000000_010110110;
		Dplus[942] = 18'b000000000_010110110;
		Dplus[943] = 18'b000000000_010110110;
		Dplus[944] = 18'b000000000_010110110;
		Dplus[945] = 18'b000000000_010110101;
		Dplus[946] = 18'b000000000_010110101;
		Dplus[947] = 18'b000000000_010110101;
		Dplus[948] = 18'b000000000_010110101;
		Dplus[949] = 18'b000000000_010110100;
		Dplus[950] = 18'b000000000_010110100;
		Dplus[951] = 18'b000000000_010110100;
		Dplus[952] = 18'b000000000_010110100;
		Dplus[953] = 18'b000000000_010110100;
		Dplus[954] = 18'b000000000_010110011;
		Dplus[955] = 18'b000000000_010110011;
		Dplus[956] = 18'b000000000_010110011;
		Dplus[957] = 18'b000000000_010110011;
		Dplus[958] = 18'b000000000_010110011;
		Dplus[959] = 18'b000000000_010110010;
		Dplus[960] = 18'b000000000_010110010;
		Dplus[961] = 18'b000000000_010110010;
		Dplus[962] = 18'b000000000_010110010;
		Dplus[963] = 18'b000000000_010110001;
		Dplus[964] = 18'b000000000_010110001;
		Dplus[965] = 18'b000000000_010110001;
		Dplus[966] = 18'b000000000_010110001;
		Dplus[967] = 18'b000000000_010110001;
		Dplus[968] = 18'b000000000_010110000;
		Dplus[969] = 18'b000000000_010110000;
		Dplus[970] = 18'b000000000_010110000;
		Dplus[971] = 18'b000000000_010110000;
		Dplus[972] = 18'b000000000_010110000;
		Dplus[973] = 18'b000000000_010101111;
		Dplus[974] = 18'b000000000_010101111;
		Dplus[975] = 18'b000000000_010101111;
		Dplus[976] = 18'b000000000_010101111;
		Dplus[977] = 18'b000000000_010101110;
		Dplus[978] = 18'b000000000_010101110;
		Dplus[979] = 18'b000000000_010101110;
		Dplus[980] = 18'b000000000_010101110;
		Dplus[981] = 18'b000000000_010101110;
		Dplus[982] = 18'b000000000_010101101;
		Dplus[983] = 18'b000000000_010101101;
		Dplus[984] = 18'b000000000_010101101;
		Dplus[985] = 18'b000000000_010101101;
		Dplus[986] = 18'b000000000_010101101;
		Dplus[987] = 18'b000000000_010101100;
		Dplus[988] = 18'b000000000_010101100;
		Dplus[989] = 18'b000000000_010101100;
		Dplus[990] = 18'b000000000_010101100;
		Dplus[991] = 18'b000000000_010101100;
		Dplus[992] = 18'b000000000_010101011;
		Dplus[993] = 18'b000000000_010101011;
		Dplus[994] = 18'b000000000_010101011;
		Dplus[995] = 18'b000000000_010101011;
		Dplus[996] = 18'b000000000_010101011;
		Dplus[997] = 18'b000000000_010101010;
		Dplus[998] = 18'b000000000_010101010;
		Dplus[999] = 18'b000000000_010101010;
		Dplus[1000] = 18'b000000000_010101010;
		Dplus[1001] = 18'b000000000_010101001;
		Dplus[1002] = 18'b000000000_010101001;
		Dplus[1003] = 18'b000000000_010101001;
		Dplus[1004] = 18'b000000000_010101001;
		Dplus[1005] = 18'b000000000_010101001;
		Dplus[1006] = 18'b000000000_010101000;
		Dplus[1007] = 18'b000000000_010101000;
		Dplus[1008] = 18'b000000000_010101000;
		Dplus[1009] = 18'b000000000_010101000;
		Dplus[1010] = 18'b000000000_010101000;
		Dplus[1011] = 18'b000000000_010100111;
		Dplus[1012] = 18'b000000000_010100111;
		Dplus[1013] = 18'b000000000_010100111;
		Dplus[1014] = 18'b000000000_010100111;
		Dplus[1015] = 18'b000000000_010100111;
		Dplus[1016] = 18'b000000000_010100110;
		Dplus[1017] = 18'b000000000_010100110;
		Dplus[1018] = 18'b000000000_010100110;
		Dplus[1019] = 18'b000000000_010100110;
		Dplus[1020] = 18'b000000000_010100110;
		Dplus[1021] = 18'b000000000_010100101;
		Dplus[1022] = 18'b000000000_010100101;
		Dplus[1023] = 18'b000000000_010100101;
		DplusInteger[2] = 18'b000000000_010100101;
		DplusInteger[3] = 18'b000000000_001010111;
		DplusInteger[4] = 18'b000000000_000101101;
		DplusInteger[5] = 18'b000000000_000010111;
		DplusInteger[6] = 18'b000000000_000001011;
		DplusInteger[7] = 18'b000000000_000000110;
		DplusInteger[8] = 18'b000000000_000000011;
		DplusInteger[9] = 18'b000000000_000000001;
		DplusInteger[10] = 18'b000000000_000000001;
		DplusInteger[11] = 18'b000000000_000000000;
		DplusInteger[12] = 18'b000000000_000000000;
		DplusInteger[13] = 18'b000000000_000000000;
		DplusInteger[14] = 18'b000000000_000000000;
		DplusInteger[15] = 18'b000000000_000000000;
		DplusInteger[16] = 18'b000000000_000000000;
		DplusInteger[17] = 18'b000000000_000000000;
		DplusInteger[18] = 18'b000000000_000000000;
		DplusInteger[19] = 18'b000000000_000000000;
		DplusInteger[20] = 18'b000000000_000000000;
		DplusInteger[21] = 18'b000000000_000000000;
		DplusInteger[22] = 18'b000000000_000000000;
		DplusInteger[23] = 18'b000000000_000000000;
		DplusInteger[24] = 18'b000000000_000000000;
		DplusInteger[25] = 18'b000000000_000000000;
		DplusInteger[26] = 18'b000000000_000000000;
		DplusInteger[27] = 18'b000000000_000000000;
		DplusInteger[28] = 18'b000000000_000000000;
		DplusInteger[29] = 18'b000000000_000000000;
		DplusInteger[30] = 18'b000000000_000000000;
		DplusInteger[31] = 18'b000000000_000000000;
		DplusInteger[32] = 18'b000000000_000000000;
		DplusInteger[33] = 18'b000000000_000000000;
		DplusInteger[34] = 18'b000000000_000000000;
		DplusInteger[35] = 18'b000000000_000000000;
		DplusInteger[36] = 18'b000000000_000000000;
		DplusInteger[37] = 18'b000000000_000000000;
		DplusInteger[38] = 18'b000000000_000000000;
		DplusInteger[39] = 18'b000000000_000000000;
		DplusInteger[40] = 18'b000000000_000000000;
		DplusInteger[41] = 18'b000000000_000000000;
		DplusInteger[42] = 18'b000000000_000000000;
		DplusInteger[43] = 18'b000000000_000000000;
		DplusInteger[44] = 18'b000000000_000000000;
		DplusInteger[45] = 18'b000000000_000000000;
		DplusInteger[46] = 18'b000000000_000000000;
		DplusInteger[47] = 18'b000000000_000000000;
		DplusInteger[48] = 18'b000000000_000000000;
		DplusInteger[49] = 18'b000000000_000000000;
		DplusInteger[50] = 18'b000000000_000000000;
		DplusInteger[51] = 18'b000000000_000000000;
		DplusInteger[52] = 18'b000000000_000000000;
		DplusInteger[53] = 18'b000000000_000000000;
		DplusInteger[54] = 18'b000000000_000000000;
		DplusInteger[55] = 18'b000000000_000000000;
		DplusInteger[56] = 18'b000000000_000000000;
		DplusInteger[57] = 18'b000000000_000000000;
		DplusInteger[58] = 18'b000000000_000000000;
		DplusInteger[59] = 18'b000000000_000000000;
		DplusInteger[60] = 18'b000000000_000000000;
		DplusInteger[61] = 18'b000000000_000000000;
		DplusInteger[62] = 18'b000000000_000000000;
		DplusInteger[63] = 18'b000000000_000000000;
		DplusInteger[64] = 18'b000000000_000000000;
		DplusInteger[65] = 18'b000000000_000000000;
		DplusInteger[66] = 18'b000000000_000000000;
		DplusInteger[67] = 18'b000000000_000000000;
		DplusInteger[68] = 18'b000000000_000000000;
		DplusInteger[69] = 18'b000000000_000000000;
		DplusInteger[70] = 18'b000000000_000000000;
		DplusInteger[71] = 18'b000000000_000000000;
		DplusInteger[72] = 18'b000000000_000000000;
		DplusInteger[73] = 18'b000000000_000000000;
		DplusInteger[74] = 18'b000000000_000000000;
		DplusInteger[75] = 18'b000000000_000000000;
		DplusInteger[76] = 18'b000000000_000000000;
		DplusInteger[77] = 18'b000000000_000000000;
		DplusInteger[78] = 18'b000000000_000000000;
		DplusInteger[79] = 18'b000000000_000000000;
		DplusInteger[80] = 18'b000000000_000000000;
		DplusInteger[81] = 18'b000000000_000000000;
		DplusInteger[82] = 18'b000000000_000000000;
		DplusInteger[83] = 18'b000000000_000000000;
		DplusInteger[84] = 18'b000000000_000000000;
		DplusInteger[85] = 18'b000000000_000000000;
		DplusInteger[86] = 18'b000000000_000000000;
		DplusInteger[87] = 18'b000000000_000000000;
		DplusInteger[88] = 18'b000000000_000000000;
		DplusInteger[89] = 18'b000000000_000000000;
		DplusInteger[90] = 18'b000000000_000000000;
		DplusInteger[91] = 18'b000000000_000000000;
		DplusInteger[92] = 18'b000000000_000000000;
		DplusInteger[93] = 18'b000000000_000000000;
		DplusInteger[94] = 18'b000000000_000000000;
		DplusInteger[95] = 18'b000000000_000000000;
		DplusInteger[96] = 18'b000000000_000000000;
		DplusInteger[97] = 18'b000000000_000000000;
		DplusInteger[98] = 18'b000000000_000000000;
		DplusInteger[99] = 18'b000000000_000000000;
		DplusInteger[100] = 18'b000000000_000000000;
		DplusInteger[101] = 18'b000000000_000000000;
		DplusInteger[102] = 18'b000000000_000000000;
		DplusInteger[103] = 18'b000000000_000000000;
		DplusInteger[104] = 18'b000000000_000000000;
		DplusInteger[105] = 18'b000000000_000000000;
		DplusInteger[106] = 18'b000000000_000000000;
		DplusInteger[107] = 18'b000000000_000000000;
		DplusInteger[108] = 18'b000000000_000000000;
		DplusInteger[109] = 18'b000000000_000000000;
		DplusInteger[110] = 18'b000000000_000000000;
		DplusInteger[111] = 18'b000000000_000000000;
		DplusInteger[112] = 18'b000000000_000000000;
		DplusInteger[113] = 18'b000000000_000000000;
		DplusInteger[114] = 18'b000000000_000000000;
		DplusInteger[115] = 18'b000000000_000000000;
		DplusInteger[116] = 18'b000000000_000000000;
		DplusInteger[117] = 18'b000000000_000000000;
		DplusInteger[118] = 18'b000000000_000000000;
		DplusInteger[119] = 18'b000000000_000000000;
		DplusInteger[120] = 18'b000000000_000000000;
		DplusInteger[121] = 18'b000000000_000000000;
		DplusInteger[122] = 18'b000000000_000000000;
		DplusInteger[123] = 18'b000000000_000000000;
		DplusInteger[124] = 18'b000000000_000000000;
		DplusInteger[125] = 18'b000000000_000000000;
		DplusInteger[126] = 18'b000000000_000000000;
		DplusInteger[127] = 18'b000000000_000000000;
		DplusInteger[128] = 18'b000000000_000000000;
		DplusInteger[129] = 18'b000000000_000000000;
		DplusInteger[130] = 18'b000000000_000000000;
		DplusInteger[131] = 18'b000000000_000000000;
		DplusInteger[132] = 18'b000000000_000000000;
		DplusInteger[133] = 18'b000000000_000000000;
		DplusInteger[134] = 18'b000000000_000000000;
		DplusInteger[135] = 18'b000000000_000000000;
		DplusInteger[136] = 18'b000000000_000000000;
		DplusInteger[137] = 18'b000000000_000000000;
		DplusInteger[138] = 18'b000000000_000000000;
		DplusInteger[139] = 18'b000000000_000000000;
		DplusInteger[140] = 18'b000000000_000000000;
		DplusInteger[141] = 18'b000000000_000000000;
		DplusInteger[142] = 18'b000000000_000000000;
		DplusInteger[143] = 18'b000000000_000000000;
		DplusInteger[144] = 18'b000000000_000000000;
		DplusInteger[145] = 18'b000000000_000000000;
		DplusInteger[146] = 18'b000000000_000000000;
		DplusInteger[147] = 18'b000000000_000000000;
		DplusInteger[148] = 18'b000000000_000000000;
		DplusInteger[149] = 18'b000000000_000000000;
		DplusInteger[150] = 18'b000000000_000000000;
		DplusInteger[151] = 18'b000000000_000000000;
		DplusInteger[152] = 18'b000000000_000000000;
		DplusInteger[153] = 18'b000000000_000000000;
		DplusInteger[154] = 18'b000000000_000000000;
		DplusInteger[155] = 18'b000000000_000000000;
		DplusInteger[156] = 18'b000000000_000000000;
		DplusInteger[157] = 18'b000000000_000000000;
		DplusInteger[158] = 18'b000000000_000000000;
		DplusInteger[159] = 18'b000000000_000000000;
		DplusInteger[160] = 18'b000000000_000000000;
		DplusInteger[161] = 18'b000000000_000000000;
		DplusInteger[162] = 18'b000000000_000000000;
		DplusInteger[163] = 18'b000000000_000000000;
		DplusInteger[164] = 18'b000000000_000000000;
		DplusInteger[165] = 18'b000000000_000000000;
		DplusInteger[166] = 18'b000000000_000000000;
		DplusInteger[167] = 18'b000000000_000000000;
		DplusInteger[168] = 18'b000000000_000000000;
		DplusInteger[169] = 18'b000000000_000000000;
		DplusInteger[170] = 18'b000000000_000000000;
		DplusInteger[171] = 18'b000000000_000000000;
		DplusInteger[172] = 18'b000000000_000000000;
		DplusInteger[173] = 18'b000000000_000000000;
		DplusInteger[174] = 18'b000000000_000000000;
		DplusInteger[175] = 18'b000000000_000000000;
		DplusInteger[176] = 18'b000000000_000000000;
		DplusInteger[177] = 18'b000000000_000000000;
		DplusInteger[178] = 18'b000000000_000000000;
		DplusInteger[179] = 18'b000000000_000000000;
		DplusInteger[180] = 18'b000000000_000000000;
		DplusInteger[181] = 18'b000000000_000000000;
		DplusInteger[182] = 18'b000000000_000000000;
		DplusInteger[183] = 18'b000000000_000000000;
		DplusInteger[184] = 18'b000000000_000000000;
		DplusInteger[185] = 18'b000000000_000000000;
		DplusInteger[186] = 18'b000000000_000000000;
		DplusInteger[187] = 18'b000000000_000000000;
		DplusInteger[188] = 18'b000000000_000000000;
		DplusInteger[189] = 18'b000000000_000000000;
		DplusInteger[190] = 18'b000000000_000000000;
		DplusInteger[191] = 18'b000000000_000000000;
		DplusInteger[192] = 18'b000000000_000000000;
		DplusInteger[193] = 18'b000000000_000000000;
		DplusInteger[194] = 18'b000000000_000000000;
		DplusInteger[195] = 18'b000000000_000000000;
		DplusInteger[196] = 18'b000000000_000000000;
		DplusInteger[197] = 18'b000000000_000000000;
		DplusInteger[198] = 18'b000000000_000000000;
		DplusInteger[199] = 18'b000000000_000000000;
		DplusInteger[200] = 18'b000000000_000000000;
		DplusInteger[201] = 18'b000000000_000000000;
		DplusInteger[202] = 18'b000000000_000000000;
		DplusInteger[203] = 18'b000000000_000000000;
		DplusInteger[204] = 18'b000000000_000000000;
		DplusInteger[205] = 18'b000000000_000000000;
		DplusInteger[206] = 18'b000000000_000000000;
		DplusInteger[207] = 18'b000000000_000000000;
		DplusInteger[208] = 18'b000000000_000000000;
		DplusInteger[209] = 18'b000000000_000000000;
		DplusInteger[210] = 18'b000000000_000000000;
		DplusInteger[211] = 18'b000000000_000000000;
		DplusInteger[212] = 18'b000000000_000000000;
		DplusInteger[213] = 18'b000000000_000000000;
		DplusInteger[214] = 18'b000000000_000000000;
		DplusInteger[215] = 18'b000000000_000000000;
		DplusInteger[216] = 18'b000000000_000000000;
		DplusInteger[217] = 18'b000000000_000000000;
		DplusInteger[218] = 18'b000000000_000000000;
		DplusInteger[219] = 18'b000000000_000000000;
		DplusInteger[220] = 18'b000000000_000000000;
		DplusInteger[221] = 18'b000000000_000000000;
		DplusInteger[222] = 18'b000000000_000000000;
		DplusInteger[223] = 18'b000000000_000000000;
		DplusInteger[224] = 18'b000000000_000000000;
		DplusInteger[225] = 18'b000000000_000000000;
		DplusInteger[226] = 18'b000000000_000000000;
		DplusInteger[227] = 18'b000000000_000000000;
		DplusInteger[228] = 18'b000000000_000000000;
		DplusInteger[229] = 18'b000000000_000000000;
		DplusInteger[230] = 18'b000000000_000000000;
		DplusInteger[231] = 18'b000000000_000000000;
		DplusInteger[232] = 18'b000000000_000000000;
		DplusInteger[233] = 18'b000000000_000000000;
		DplusInteger[234] = 18'b000000000_000000000;
		DplusInteger[235] = 18'b000000000_000000000;
		DplusInteger[236] = 18'b000000000_000000000;
		DplusInteger[237] = 18'b000000000_000000000;
		DplusInteger[238] = 18'b000000000_000000000;
		DplusInteger[239] = 18'b000000000_000000000;
		DplusInteger[240] = 18'b000000000_000000000;
		DplusInteger[241] = 18'b000000000_000000000;
		DplusInteger[242] = 18'b000000000_000000000;
		DplusInteger[243] = 18'b000000000_000000000;
		DplusInteger[244] = 18'b000000000_000000000;
		DplusInteger[245] = 18'b000000000_000000000;
		DplusInteger[246] = 18'b000000000_000000000;
		DplusInteger[247] = 18'b000000000_000000000;
		DplusInteger[248] = 18'b000000000_000000000;
		DplusInteger[249] = 18'b000000000_000000000;
		DplusInteger[250] = 18'b000000000_000000000;
		DplusInteger[251] = 18'b000000000_000000000;
		DplusInteger[252] = 18'b000000000_000000000;
		DplusInteger[253] = 18'b000000000_000000000;
		DplusInteger[254] = 18'b000000000_000000000;
		DplusInteger[255] = 18'b000000000_000000000;
		DminusInteger[2] = 18'b111111111_100101100;
		DminusInteger[3] = 18'b111111111_110011101;
		DminusInteger[4] = 18'b111111111_111010000;
		DminusInteger[5] = 18'b111111111_111101001;
		DminusInteger[6] = 18'b111111111_111110100;
		DminusInteger[7] = 18'b111111111_111111010;
		DminusInteger[8] = 18'b111111111_111111101;
		DminusInteger[9] = 18'b111111111_111111111;
		DminusInteger[10] = 18'b111111111_111111111;
		DminusInteger[11] = 18'b000000000_000000000;
		DminusInteger[12] = 18'b000000000_000000000;
		DminusInteger[13] = 18'b000000000_000000000;
		DminusInteger[14] = 18'b000000000_000000000;
		DminusInteger[15] = 18'b000000000_000000000;
		DminusInteger[16] = 18'b000000000_000000000;
		DminusInteger[17] = 18'b000000000_000000000;
		DminusInteger[18] = 18'b000000000_000000000;
		DminusInteger[19] = 18'b000000000_000000000;
		DminusInteger[20] = 18'b000000000_000000000;
		DminusInteger[21] = 18'b000000000_000000000;
		DminusInteger[22] = 18'b000000000_000000000;
		DminusInteger[23] = 18'b000000000_000000000;
		DminusInteger[24] = 18'b000000000_000000000;
		DminusInteger[25] = 18'b000000000_000000000;
		DminusInteger[26] = 18'b000000000_000000000;
		DminusInteger[27] = 18'b000000000_000000000;
		DminusInteger[28] = 18'b000000000_000000000;
		DminusInteger[29] = 18'b000000000_000000000;
		DminusInteger[30] = 18'b000000000_000000000;
		DminusInteger[31] = 18'b000000000_000000000;
		DminusInteger[32] = 18'b000000000_000000000;
		DminusInteger[33] = 18'b000000000_000000000;
		DminusInteger[34] = 18'b000000000_000000000;
		DminusInteger[35] = 18'b000000000_000000000;
		DminusInteger[36] = 18'b000000000_000000000;
		DminusInteger[37] = 18'b000000000_000000000;
		DminusInteger[38] = 18'b000000000_000000000;
		DminusInteger[39] = 18'b000000000_000000000;
		DminusInteger[40] = 18'b000000000_000000000;
		DminusInteger[41] = 18'b000000000_000000000;
		DminusInteger[42] = 18'b000000000_000000000;
		DminusInteger[43] = 18'b000000000_000000000;
		DminusInteger[44] = 18'b000000000_000000000;
		DminusInteger[45] = 18'b000000000_000000000;
		DminusInteger[46] = 18'b000000000_000000000;
		DminusInteger[47] = 18'b000000000_000000000;
		DminusInteger[48] = 18'b000000000_000000000;
		DminusInteger[49] = 18'b000000000_000000000;
		DminusInteger[50] = 18'b000000000_000000000;
		DminusInteger[51] = 18'b000000000_000000000;
		DminusInteger[52] = 18'b000000000_000000000;
		DminusInteger[53] = 18'b000000000_000000000;
		DminusInteger[54] = 18'b000000000_000000000;
		DminusInteger[55] = 18'b000000000_000000000;
		DminusInteger[56] = 18'b000000000_000000000;
		DminusInteger[57] = 18'b000000000_000000000;
		DminusInteger[58] = 18'b000000000_000000000;
		DminusInteger[59] = 18'b000000000_000000000;
		DminusInteger[60] = 18'b000000000_000000000;
		DminusInteger[61] = 18'b000000000_000000000;
		DminusInteger[62] = 18'b000000000_000000000;
		DminusInteger[63] = 18'b000000000_000000000;
		DminusInteger[64] = 18'b000000000_000000000;
		DminusInteger[65] = 18'b000000000_000000000;
		DminusInteger[66] = 18'b000000000_000000000;
		DminusInteger[67] = 18'b000000000_000000000;
		DminusInteger[68] = 18'b000000000_000000000;
		DminusInteger[69] = 18'b000000000_000000000;
		DminusInteger[70] = 18'b000000000_000000000;
		DminusInteger[71] = 18'b000000000_000000000;
		DminusInteger[72] = 18'b000000000_000000000;
		DminusInteger[73] = 18'b000000000_000000000;
		DminusInteger[74] = 18'b000000000_000000000;
		DminusInteger[75] = 18'b000000000_000000000;
		DminusInteger[76] = 18'b000000000_000000000;
		DminusInteger[77] = 18'b000000000_000000000;
		DminusInteger[78] = 18'b000000000_000000000;
		DminusInteger[79] = 18'b000000000_000000000;
		DminusInteger[80] = 18'b000000000_000000000;
		DminusInteger[81] = 18'b000000000_000000000;
		DminusInteger[82] = 18'b000000000_000000000;
		DminusInteger[83] = 18'b000000000_000000000;
		DminusInteger[84] = 18'b000000000_000000000;
		DminusInteger[85] = 18'b000000000_000000000;
		DminusInteger[86] = 18'b000000000_000000000;
		DminusInteger[87] = 18'b000000000_000000000;
		DminusInteger[88] = 18'b000000000_000000000;
		DminusInteger[89] = 18'b000000000_000000000;
		DminusInteger[90] = 18'b000000000_000000000;
		DminusInteger[91] = 18'b000000000_000000000;
		DminusInteger[92] = 18'b000000000_000000000;
		DminusInteger[93] = 18'b000000000_000000000;
		DminusInteger[94] = 18'b000000000_000000000;
		DminusInteger[95] = 18'b000000000_000000000;
		DminusInteger[96] = 18'b000000000_000000000;
		DminusInteger[97] = 18'b000000000_000000000;
		DminusInteger[98] = 18'b000000000_000000000;
		DminusInteger[99] = 18'b000000000_000000000;
		DminusInteger[100] = 18'b000000000_000000000;
		DminusInteger[101] = 18'b000000000_000000000;
		DminusInteger[102] = 18'b000000000_000000000;
		DminusInteger[103] = 18'b000000000_000000000;
		DminusInteger[104] = 18'b000000000_000000000;
		DminusInteger[105] = 18'b000000000_000000000;
		DminusInteger[106] = 18'b000000000_000000000;
		DminusInteger[107] = 18'b000000000_000000000;
		DminusInteger[108] = 18'b000000000_000000000;
		DminusInteger[109] = 18'b000000000_000000000;
		DminusInteger[110] = 18'b000000000_000000000;
		DminusInteger[111] = 18'b000000000_000000000;
		DminusInteger[112] = 18'b000000000_000000000;
		DminusInteger[113] = 18'b000000000_000000000;
		DminusInteger[114] = 18'b000000000_000000000;
		DminusInteger[115] = 18'b000000000_000000000;
		DminusInteger[116] = 18'b000000000_000000000;
		DminusInteger[117] = 18'b000000000_000000000;
		DminusInteger[118] = 18'b000000000_000000000;
		DminusInteger[119] = 18'b000000000_000000000;
		DminusInteger[120] = 18'b000000000_000000000;
		DminusInteger[121] = 18'b000000000_000000000;
		DminusInteger[122] = 18'b000000000_000000000;
		DminusInteger[123] = 18'b000000000_000000000;
		DminusInteger[124] = 18'b000000000_000000000;
		DminusInteger[125] = 18'b000000000_000000000;
		DminusInteger[126] = 18'b000000000_000000000;
		DminusInteger[127] = 18'b000000000_000000000;
		DminusInteger[128] = 18'b000000000_000000000;
		DminusInteger[129] = 18'b000000000_000000000;
		DminusInteger[130] = 18'b000000000_000000000;
		DminusInteger[131] = 18'b000000000_000000000;
		DminusInteger[132] = 18'b000000000_000000000;
		DminusInteger[133] = 18'b000000000_000000000;
		DminusInteger[134] = 18'b000000000_000000000;
		DminusInteger[135] = 18'b000000000_000000000;
		DminusInteger[136] = 18'b000000000_000000000;
		DminusInteger[137] = 18'b000000000_000000000;
		DminusInteger[138] = 18'b000000000_000000000;
		DminusInteger[139] = 18'b000000000_000000000;
		DminusInteger[140] = 18'b000000000_000000000;
		DminusInteger[141] = 18'b000000000_000000000;
		DminusInteger[142] = 18'b000000000_000000000;
		DminusInteger[143] = 18'b000000000_000000000;
		DminusInteger[144] = 18'b000000000_000000000;
		DminusInteger[145] = 18'b000000000_000000000;
		DminusInteger[146] = 18'b000000000_000000000;
		DminusInteger[147] = 18'b000000000_000000000;
		DminusInteger[148] = 18'b000000000_000000000;
		DminusInteger[149] = 18'b000000000_000000000;
		DminusInteger[150] = 18'b000000000_000000000;
		DminusInteger[151] = 18'b000000000_000000000;
		DminusInteger[152] = 18'b000000000_000000000;
		DminusInteger[153] = 18'b000000000_000000000;
		DminusInteger[154] = 18'b000000000_000000000;
		DminusInteger[155] = 18'b000000000_000000000;
		DminusInteger[156] = 18'b000000000_000000000;
		DminusInteger[157] = 18'b000000000_000000000;
		DminusInteger[158] = 18'b000000000_000000000;
		DminusInteger[159] = 18'b000000000_000000000;
		DminusInteger[160] = 18'b000000000_000000000;
		DminusInteger[161] = 18'b000000000_000000000;
		DminusInteger[162] = 18'b000000000_000000000;
		DminusInteger[163] = 18'b000000000_000000000;
		DminusInteger[164] = 18'b000000000_000000000;
		DminusInteger[165] = 18'b000000000_000000000;
		DminusInteger[166] = 18'b000000000_000000000;
		DminusInteger[167] = 18'b000000000_000000000;
		DminusInteger[168] = 18'b000000000_000000000;
		DminusInteger[169] = 18'b000000000_000000000;
		DminusInteger[170] = 18'b000000000_000000000;
		DminusInteger[171] = 18'b000000000_000000000;
		DminusInteger[172] = 18'b000000000_000000000;
		DminusInteger[173] = 18'b000000000_000000000;
		DminusInteger[174] = 18'b000000000_000000000;
		DminusInteger[175] = 18'b000000000_000000000;
		DminusInteger[176] = 18'b000000000_000000000;
		DminusInteger[177] = 18'b000000000_000000000;
		DminusInteger[178] = 18'b000000000_000000000;
		DminusInteger[179] = 18'b000000000_000000000;
		DminusInteger[180] = 18'b000000000_000000000;
		DminusInteger[181] = 18'b000000000_000000000;
		DminusInteger[182] = 18'b000000000_000000000;
		DminusInteger[183] = 18'b000000000_000000000;
		DminusInteger[184] = 18'b000000000_000000000;
		DminusInteger[185] = 18'b000000000_000000000;
		DminusInteger[186] = 18'b000000000_000000000;
		DminusInteger[187] = 18'b000000000_000000000;
		DminusInteger[188] = 18'b000000000_000000000;
		DminusInteger[189] = 18'b000000000_000000000;
		DminusInteger[190] = 18'b000000000_000000000;
		DminusInteger[191] = 18'b000000000_000000000;
		DminusInteger[192] = 18'b000000000_000000000;
		DminusInteger[193] = 18'b000000000_000000000;
		DminusInteger[194] = 18'b000000000_000000000;
		DminusInteger[195] = 18'b000000000_000000000;
		DminusInteger[196] = 18'b000000000_000000000;
		DminusInteger[197] = 18'b000000000_000000000;
		DminusInteger[198] = 18'b000000000_000000000;
		DminusInteger[199] = 18'b000000000_000000000;
		DminusInteger[200] = 18'b000000000_000000000;
		DminusInteger[201] = 18'b000000000_000000000;
		DminusInteger[202] = 18'b000000000_000000000;
		DminusInteger[203] = 18'b000000000_000000000;
		DminusInteger[204] = 18'b000000000_000000000;
		DminusInteger[205] = 18'b000000000_000000000;
		DminusInteger[206] = 18'b000000000_000000000;
		DminusInteger[207] = 18'b000000000_000000000;
		DminusInteger[208] = 18'b000000000_000000000;
		DminusInteger[209] = 18'b000000000_000000000;
		DminusInteger[210] = 18'b000000000_000000000;
		DminusInteger[211] = 18'b000000000_000000000;
		DminusInteger[212] = 18'b000000000_000000000;
		DminusInteger[213] = 18'b000000000_000000000;
		DminusInteger[214] = 18'b000000000_000000000;
		DminusInteger[215] = 18'b000000000_000000000;
		DminusInteger[216] = 18'b000000000_000000000;
		DminusInteger[217] = 18'b000000000_000000000;
		DminusInteger[218] = 18'b000000000_000000000;
		DminusInteger[219] = 18'b000000000_000000000;
		DminusInteger[220] = 18'b000000000_000000000;
		DminusInteger[221] = 18'b000000000_000000000;
		DminusInteger[222] = 18'b000000000_000000000;
		DminusInteger[223] = 18'b000000000_000000000;
		DminusInteger[224] = 18'b000000000_000000000;
		DminusInteger[225] = 18'b000000000_000000000;
		DminusInteger[226] = 18'b000000000_000000000;
		DminusInteger[227] = 18'b000000000_000000000;
		DminusInteger[228] = 18'b000000000_000000000;
		DminusInteger[229] = 18'b000000000_000000000;
		DminusInteger[230] = 18'b000000000_000000000;
		DminusInteger[231] = 18'b000000000_000000000;
		DminusInteger[232] = 18'b000000000_000000000;
		DminusInteger[233] = 18'b000000000_000000000;
		DminusInteger[234] = 18'b000000000_000000000;
		DminusInteger[235] = 18'b000000000_000000000;
		DminusInteger[236] = 18'b000000000_000000000;
		DminusInteger[237] = 18'b000000000_000000000;
		DminusInteger[238] = 18'b000000000_000000000;
		DminusInteger[239] = 18'b000000000_000000000;
		DminusInteger[240] = 18'b000000000_000000000;
		DminusInteger[241] = 18'b000000000_000000000;
		DminusInteger[242] = 18'b000000000_000000000;
		DminusInteger[243] = 18'b000000000_000000000;
		DminusInteger[244] = 18'b000000000_000000000;
		DminusInteger[245] = 18'b000000000_000000000;
		DminusInteger[246] = 18'b000000000_000000000;
		DminusInteger[247] = 18'b000000000_000000000;
		DminusInteger[248] = 18'b000000000_000000000;
		DminusInteger[249] = 18'b000000000_000000000;
		DminusInteger[250] = 18'b000000000_000000000;
		DminusInteger[251] = 18'b000000000_000000000;
		DminusInteger[252] = 18'b000000000_000000000;
		DminusInteger[253] = 18'b000000000_000000000;
		DminusInteger[254] = 18'b000000000_000000000;
		DminusInteger[255] = 18'b000000000_000000000;
end
endmodule
