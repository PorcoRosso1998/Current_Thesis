module Tables();
	reg [15:0] Dplus[511:0];
	reg [15:0] Dminus[511:0];
	reg [7:0] DminusInteger[127:0];
	reg [7:0] DplusInteger[127:0];
	initial begin
		Dminus[1] = 16'b11110111_01111000;
		Dminus[2] = 16'b11111000_01111000;
		Dminus[3] = 16'b11111001_00001101;
		Dminus[4] = 16'b11111001_01110111;
		Dminus[5] = 16'b11111001_11001001;
		Dminus[6] = 16'b11111010_00001011;
		Dminus[7] = 16'b11111010_01000100;
		Dminus[8] = 16'b11111010_01110101;
		Dminus[9] = 16'b11111010_10100000;
		Dminus[10] = 16'b11111010_11000110;
		Dminus[11] = 16'b11111010_11101001;
		Dminus[12] = 16'b11111011_00001000;
		Dminus[13] = 16'b11111011_00100101;
		Dminus[14] = 16'b11111011_01000000;
		Dminus[15] = 16'b11111011_01011001;
		Dminus[16] = 16'b11111011_01110001;
		Dminus[17] = 16'b11111011_10000111;
		Dminus[18] = 16'b11111011_10011011;
		Dminus[19] = 16'b11111011_10101111;
		Dminus[20] = 16'b11111011_11000001;
		Dminus[21] = 16'b11111011_11010011;
		Dminus[22] = 16'b11111011_11100011;
		Dminus[23] = 16'b11111011_11110011;
		Dminus[24] = 16'b11111100_00000010;
		Dminus[25] = 16'b11111100_00010001;
		Dminus[26] = 16'b11111100_00011111;
		Dminus[27] = 16'b11111100_00101100;
		Dminus[28] = 16'b11111100_00111001;
		Dminus[29] = 16'b11111100_01000110;
		Dminus[30] = 16'b11111100_01010010;
		Dminus[31] = 16'b11111100_01011110;
		Dminus[32] = 16'b11111100_01101001;
		Dminus[33] = 16'b11111100_01110100;
		Dminus[34] = 16'b11111100_01111110;
		Dminus[35] = 16'b11111100_10001000;
		Dminus[36] = 16'b11111100_10010010;
		Dminus[37] = 16'b11111100_10011100;
		Dminus[38] = 16'b11111100_10100101;
		Dminus[39] = 16'b11111100_10101110;
		Dminus[40] = 16'b11111100_10110111;
		Dminus[41] = 16'b11111100_11000000;
		Dminus[42] = 16'b11111100_11001000;
		Dminus[43] = 16'b11111100_11010000;
		Dminus[44] = 16'b11111100_11011000;
		Dminus[45] = 16'b11111100_11100000;
		Dminus[46] = 16'b11111100_11101000;
		Dminus[47] = 16'b11111100_11101111;
		Dminus[48] = 16'b11111100_11110111;
		Dminus[49] = 16'b11111100_11111110;
		Dminus[50] = 16'b11111101_00000101;
		Dminus[51] = 16'b11111101_00001100;
		Dminus[52] = 16'b11111101_00010010;
		Dminus[53] = 16'b11111101_00011001;
		Dminus[54] = 16'b11111101_00011111;
		Dminus[55] = 16'b11111101_00100110;
		Dminus[56] = 16'b11111101_00101100;
		Dminus[57] = 16'b11111101_00110010;
		Dminus[58] = 16'b11111101_00111000;
		Dminus[59] = 16'b11111101_00111101;
		Dminus[60] = 16'b11111101_01000011;
		Dminus[61] = 16'b11111101_01001001;
		Dminus[62] = 16'b11111101_01001110;
		Dminus[63] = 16'b11111101_01010100;
		Dminus[64] = 16'b11111101_01011001;
		Dminus[65] = 16'b11111101_01011110;
		Dminus[66] = 16'b11111101_01100011;
		Dminus[67] = 16'b11111101_01101001;
		Dminus[68] = 16'b11111101_01101110;
		Dminus[69] = 16'b11111101_01110010;
		Dminus[70] = 16'b11111101_01110111;
		Dminus[71] = 16'b11111101_01111100;
		Dminus[72] = 16'b11111101_10000001;
		Dminus[73] = 16'b11111101_10000101;
		Dminus[74] = 16'b11111101_10001010;
		Dminus[75] = 16'b11111101_10001110;
		Dminus[76] = 16'b11111101_10010011;
		Dminus[77] = 16'b11111101_10010111;
		Dminus[78] = 16'b11111101_10011011;
		Dminus[79] = 16'b11111101_10100000;
		Dminus[80] = 16'b11111101_10100100;
		Dminus[81] = 16'b11111101_10101000;
		Dminus[82] = 16'b11111101_10101100;
		Dminus[83] = 16'b11111101_10110000;
		Dminus[84] = 16'b11111101_10110100;
		Dminus[85] = 16'b11111101_10111000;
		Dminus[86] = 16'b11111101_10111100;
		Dminus[87] = 16'b11111101_10111111;
		Dminus[88] = 16'b11111101_11000011;
		Dminus[89] = 16'b11111101_11000111;
		Dminus[90] = 16'b11111101_11001010;
		Dminus[91] = 16'b11111101_11001110;
		Dminus[92] = 16'b11111101_11010010;
		Dminus[93] = 16'b11111101_11010101;
		Dminus[94] = 16'b11111101_11011001;
		Dminus[95] = 16'b11111101_11011100;
		Dminus[96] = 16'b11111101_11011111;
		Dminus[97] = 16'b11111101_11100011;
		Dminus[98] = 16'b11111101_11100110;
		Dminus[99] = 16'b11111101_11101001;
		Dminus[100] = 16'b11111101_11101101;
		Dminus[101] = 16'b11111101_11110000;
		Dminus[102] = 16'b11111101_11110011;
		Dminus[103] = 16'b11111101_11110110;
		Dminus[104] = 16'b11111101_11111001;
		Dminus[105] = 16'b11111101_11111100;
		Dminus[106] = 16'b11111101_11111111;
		Dminus[107] = 16'b11111110_00000010;
		Dminus[108] = 16'b11111110_00000101;
		Dminus[109] = 16'b11111110_00001000;
		Dminus[110] = 16'b11111110_00001011;
		Dminus[111] = 16'b11111110_00001110;
		Dminus[112] = 16'b11111110_00010001;
		Dminus[113] = 16'b11111110_00010100;
		Dminus[114] = 16'b11111110_00010110;
		Dminus[115] = 16'b11111110_00011001;
		Dminus[116] = 16'b11111110_00011100;
		Dminus[117] = 16'b11111110_00011110;
		Dminus[118] = 16'b11111110_00100001;
		Dminus[119] = 16'b11111110_00100100;
		Dminus[120] = 16'b11111110_00100110;
		Dminus[121] = 16'b11111110_00101001;
		Dminus[122] = 16'b11111110_00101100;
		Dminus[123] = 16'b11111110_00101110;
		Dminus[124] = 16'b11111110_00110001;
		Dminus[125] = 16'b11111110_00110011;
		Dminus[126] = 16'b11111110_00110110;
		Dminus[127] = 16'b11111110_00111000;
		Dminus[128] = 16'b11111110_00111010;
		Dminus[129] = 16'b11111110_00111101;
		Dminus[130] = 16'b11111110_00111111;
		Dminus[131] = 16'b11111110_01000010;
		Dminus[132] = 16'b11111110_01000100;
		Dminus[133] = 16'b11111110_01000110;
		Dminus[134] = 16'b11111110_01001001;
		Dminus[135] = 16'b11111110_01001011;
		Dminus[136] = 16'b11111110_01001101;
		Dminus[137] = 16'b11111110_01001111;
		Dminus[138] = 16'b11111110_01010010;
		Dminus[139] = 16'b11111110_01010100;
		Dminus[140] = 16'b11111110_01010110;
		Dminus[141] = 16'b11111110_01011000;
		Dminus[142] = 16'b11111110_01011010;
		Dminus[143] = 16'b11111110_01011100;
		Dminus[144] = 16'b11111110_01011110;
		Dminus[145] = 16'b11111110_01100001;
		Dminus[146] = 16'b11111110_01100011;
		Dminus[147] = 16'b11111110_01100101;
		Dminus[148] = 16'b11111110_01100111;
		Dminus[149] = 16'b11111110_01101001;
		Dminus[150] = 16'b11111110_01101011;
		Dminus[151] = 16'b11111110_01101101;
		Dminus[152] = 16'b11111110_01101111;
		Dminus[153] = 16'b11111110_01110001;
		Dminus[154] = 16'b11111110_01110011;
		Dminus[155] = 16'b11111110_01110101;
		Dminus[156] = 16'b11111110_01110110;
		Dminus[157] = 16'b11111110_01111000;
		Dminus[158] = 16'b11111110_01111010;
		Dminus[159] = 16'b11111110_01111100;
		Dminus[160] = 16'b11111110_01111110;
		Dminus[161] = 16'b11111110_10000000;
		Dminus[162] = 16'b11111110_10000010;
		Dminus[163] = 16'b11111110_10000011;
		Dminus[164] = 16'b11111110_10000101;
		Dminus[165] = 16'b11111110_10000111;
		Dminus[166] = 16'b11111110_10001001;
		Dminus[167] = 16'b11111110_10001011;
		Dminus[168] = 16'b11111110_10001100;
		Dminus[169] = 16'b11111110_10001110;
		Dminus[170] = 16'b11111110_10010000;
		Dminus[171] = 16'b11111110_10010001;
		Dminus[172] = 16'b11111110_10010011;
		Dminus[173] = 16'b11111110_10010101;
		Dminus[174] = 16'b11111110_10010110;
		Dminus[175] = 16'b11111110_10011000;
		Dminus[176] = 16'b11111110_10011010;
		Dminus[177] = 16'b11111110_10011011;
		Dminus[178] = 16'b11111110_10011101;
		Dminus[179] = 16'b11111110_10011111;
		Dminus[180] = 16'b11111110_10100000;
		Dminus[181] = 16'b11111110_10100010;
		Dminus[182] = 16'b11111110_10100011;
		Dminus[183] = 16'b11111110_10100101;
		Dminus[184] = 16'b11111110_10100110;
		Dminus[185] = 16'b11111110_10101000;
		Dminus[186] = 16'b11111110_10101010;
		Dminus[187] = 16'b11111110_10101011;
		Dminus[188] = 16'b11111110_10101101;
		Dminus[189] = 16'b11111110_10101110;
		Dminus[190] = 16'b11111110_10110000;
		Dminus[191] = 16'b11111110_10110001;
		Dminus[192] = 16'b11111110_10110011;
		Dminus[193] = 16'b11111110_10110100;
		Dminus[194] = 16'b11111110_10110101;
		Dminus[195] = 16'b11111110_10110111;
		Dminus[196] = 16'b11111110_10111000;
		Dminus[197] = 16'b11111110_10111010;
		Dminus[198] = 16'b11111110_10111011;
		Dminus[199] = 16'b11111110_10111101;
		Dminus[200] = 16'b11111110_10111110;
		Dminus[201] = 16'b11111110_10111111;
		Dminus[202] = 16'b11111110_11000001;
		Dminus[203] = 16'b11111110_11000010;
		Dminus[204] = 16'b11111110_11000011;
		Dminus[205] = 16'b11111110_11000101;
		Dminus[206] = 16'b11111110_11000110;
		Dminus[207] = 16'b11111110_11000111;
		Dminus[208] = 16'b11111110_11001001;
		Dminus[209] = 16'b11111110_11001010;
		Dminus[210] = 16'b11111110_11001011;
		Dminus[211] = 16'b11111110_11001101;
		Dminus[212] = 16'b11111110_11001110;
		Dminus[213] = 16'b11111110_11001111;
		Dminus[214] = 16'b11111110_11010001;
		Dminus[215] = 16'b11111110_11010010;
		Dminus[216] = 16'b11111110_11010011;
		Dminus[217] = 16'b11111110_11010100;
		Dminus[218] = 16'b11111110_11010110;
		Dminus[219] = 16'b11111110_11010111;
		Dminus[220] = 16'b11111110_11011000;
		Dminus[221] = 16'b11111110_11011001;
		Dminus[222] = 16'b11111110_11011011;
		Dminus[223] = 16'b11111110_11011100;
		Dminus[224] = 16'b11111110_11011101;
		Dminus[225] = 16'b11111110_11011110;
		Dminus[226] = 16'b11111110_11011111;
		Dminus[227] = 16'b11111110_11100001;
		Dminus[228] = 16'b11111110_11100010;
		Dminus[229] = 16'b11111110_11100011;
		Dminus[230] = 16'b11111110_11100100;
		Dminus[231] = 16'b11111110_11100101;
		Dminus[232] = 16'b11111110_11100110;
		Dminus[233] = 16'b11111110_11100111;
		Dminus[234] = 16'b11111110_11101001;
		Dminus[235] = 16'b11111110_11101010;
		Dminus[236] = 16'b11111110_11101011;
		Dminus[237] = 16'b11111110_11101100;
		Dminus[238] = 16'b11111110_11101101;
		Dminus[239] = 16'b11111110_11101110;
		Dminus[240] = 16'b11111110_11101111;
		Dminus[241] = 16'b11111110_11110000;
		Dminus[242] = 16'b11111110_11110001;
		Dminus[243] = 16'b11111110_11110011;
		Dminus[244] = 16'b11111110_11110100;
		Dminus[245] = 16'b11111110_11110101;
		Dminus[246] = 16'b11111110_11110110;
		Dminus[247] = 16'b11111110_11110111;
		Dminus[248] = 16'b11111110_11111000;
		Dminus[249] = 16'b11111110_11111001;
		Dminus[250] = 16'b11111110_11111010;
		Dminus[251] = 16'b11111110_11111011;
		Dminus[252] = 16'b11111110_11111100;
		Dminus[253] = 16'b11111110_11111101;
		Dminus[254] = 16'b11111110_11111110;
		Dminus[255] = 16'b11111110_11111111;
		Dminus[256] = 16'b11111111_00000000;
		Dminus[257] = 16'b11111111_00000001;
		Dminus[258] = 16'b11111111_00000010;
		Dminus[259] = 16'b11111111_00000011;
		Dminus[260] = 16'b11111111_00000100;
		Dminus[261] = 16'b11111111_00000101;
		Dminus[262] = 16'b11111111_00000110;
		Dminus[263] = 16'b11111111_00000111;
		Dminus[264] = 16'b11111111_00001000;
		Dminus[265] = 16'b11111111_00001001;
		Dminus[266] = 16'b11111111_00001010;
		Dminus[267] = 16'b11111111_00001011;
		Dminus[268] = 16'b11111111_00001100;
		Dminus[269] = 16'b11111111_00001101;
		Dminus[270] = 16'b11111111_00001101;
		Dminus[271] = 16'b11111111_00001110;
		Dminus[272] = 16'b11111111_00001111;
		Dminus[273] = 16'b11111111_00010000;
		Dminus[274] = 16'b11111111_00010001;
		Dminus[275] = 16'b11111111_00010010;
		Dminus[276] = 16'b11111111_00010011;
		Dminus[277] = 16'b11111111_00010100;
		Dminus[278] = 16'b11111111_00010101;
		Dminus[279] = 16'b11111111_00010110;
		Dminus[280] = 16'b11111111_00010111;
		Dminus[281] = 16'b11111111_00010111;
		Dminus[282] = 16'b11111111_00011000;
		Dminus[283] = 16'b11111111_00011001;
		Dminus[284] = 16'b11111111_00011010;
		Dminus[285] = 16'b11111111_00011011;
		Dminus[286] = 16'b11111111_00011100;
		Dminus[287] = 16'b11111111_00011101;
		Dminus[288] = 16'b11111111_00011101;
		Dminus[289] = 16'b11111111_00011110;
		Dminus[290] = 16'b11111111_00011111;
		Dminus[291] = 16'b11111111_00100000;
		Dminus[292] = 16'b11111111_00100001;
		Dminus[293] = 16'b11111111_00100010;
		Dminus[294] = 16'b11111111_00100010;
		Dminus[295] = 16'b11111111_00100011;
		Dminus[296] = 16'b11111111_00100100;
		Dminus[297] = 16'b11111111_00100101;
		Dminus[298] = 16'b11111111_00100110;
		Dminus[299] = 16'b11111111_00100111;
		Dminus[300] = 16'b11111111_00100111;
		Dminus[301] = 16'b11111111_00101000;
		Dminus[302] = 16'b11111111_00101001;
		Dminus[303] = 16'b11111111_00101010;
		Dminus[304] = 16'b11111111_00101010;
		Dminus[305] = 16'b11111111_00101011;
		Dminus[306] = 16'b11111111_00101100;
		Dminus[307] = 16'b11111111_00101101;
		Dminus[308] = 16'b11111111_00101110;
		Dminus[309] = 16'b11111111_00101110;
		Dminus[310] = 16'b11111111_00101111;
		Dminus[311] = 16'b11111111_00110000;
		Dminus[312] = 16'b11111111_00110001;
		Dminus[313] = 16'b11111111_00110001;
		Dminus[314] = 16'b11111111_00110010;
		Dminus[315] = 16'b11111111_00110011;
		Dminus[316] = 16'b11111111_00110100;
		Dminus[317] = 16'b11111111_00110100;
		Dminus[318] = 16'b11111111_00110101;
		Dminus[319] = 16'b11111111_00110110;
		Dminus[320] = 16'b11111111_00110111;
		Dminus[321] = 16'b11111111_00110111;
		Dminus[322] = 16'b11111111_00111000;
		Dminus[323] = 16'b11111111_00111001;
		Dminus[324] = 16'b11111111_00111001;
		Dminus[325] = 16'b11111111_00111010;
		Dminus[326] = 16'b11111111_00111011;
		Dminus[327] = 16'b11111111_00111100;
		Dminus[328] = 16'b11111111_00111100;
		Dminus[329] = 16'b11111111_00111101;
		Dminus[330] = 16'b11111111_00111110;
		Dminus[331] = 16'b11111111_00111110;
		Dminus[332] = 16'b11111111_00111111;
		Dminus[333] = 16'b11111111_01000000;
		Dminus[334] = 16'b11111111_01000000;
		Dminus[335] = 16'b11111111_01000001;
		Dminus[336] = 16'b11111111_01000010;
		Dminus[337] = 16'b11111111_01000010;
		Dminus[338] = 16'b11111111_01000011;
		Dminus[339] = 16'b11111111_01000100;
		Dminus[340] = 16'b11111111_01000100;
		Dminus[341] = 16'b11111111_01000101;
		Dminus[342] = 16'b11111111_01000110;
		Dminus[343] = 16'b11111111_01000110;
		Dminus[344] = 16'b11111111_01000111;
		Dminus[345] = 16'b11111111_01001000;
		Dminus[346] = 16'b11111111_01001000;
		Dminus[347] = 16'b11111111_01001001;
		Dminus[348] = 16'b11111111_01001010;
		Dminus[349] = 16'b11111111_01001010;
		Dminus[350] = 16'b11111111_01001011;
		Dminus[351] = 16'b11111111_01001011;
		Dminus[352] = 16'b11111111_01001100;
		Dminus[353] = 16'b11111111_01001101;
		Dminus[354] = 16'b11111111_01001101;
		Dminus[355] = 16'b11111111_01001110;
		Dminus[356] = 16'b11111111_01001111;
		Dminus[357] = 16'b11111111_01001111;
		Dminus[358] = 16'b11111111_01010000;
		Dminus[359] = 16'b11111111_01010000;
		Dminus[360] = 16'b11111111_01010001;
		Dminus[361] = 16'b11111111_01010010;
		Dminus[362] = 16'b11111111_01010010;
		Dminus[363] = 16'b11111111_01010011;
		Dminus[364] = 16'b11111111_01010011;
		Dminus[365] = 16'b11111111_01010100;
		Dminus[366] = 16'b11111111_01010101;
		Dminus[367] = 16'b11111111_01010101;
		Dminus[368] = 16'b11111111_01010110;
		Dminus[369] = 16'b11111111_01010110;
		Dminus[370] = 16'b11111111_01010111;
		Dminus[371] = 16'b11111111_01011000;
		Dminus[372] = 16'b11111111_01011000;
		Dminus[373] = 16'b11111111_01011001;
		Dminus[374] = 16'b11111111_01011001;
		Dminus[375] = 16'b11111111_01011010;
		Dminus[376] = 16'b11111111_01011010;
		Dminus[377] = 16'b11111111_01011011;
		Dminus[378] = 16'b11111111_01011100;
		Dminus[379] = 16'b11111111_01011100;
		Dminus[380] = 16'b11111111_01011101;
		Dminus[381] = 16'b11111111_01011101;
		Dminus[382] = 16'b11111111_01011110;
		Dminus[383] = 16'b11111111_01011110;
		Dminus[384] = 16'b11111111_01011111;
		Dminus[385] = 16'b11111111_01011111;
		Dminus[386] = 16'b11111111_01100000;
		Dminus[387] = 16'b11111111_01100001;
		Dminus[388] = 16'b11111111_01100001;
		Dminus[389] = 16'b11111111_01100010;
		Dminus[390] = 16'b11111111_01100010;
		Dminus[391] = 16'b11111111_01100011;
		Dminus[392] = 16'b11111111_01100011;
		Dminus[393] = 16'b11111111_01100100;
		Dminus[394] = 16'b11111111_01100100;
		Dminus[395] = 16'b11111111_01100101;
		Dminus[396] = 16'b11111111_01100101;
		Dminus[397] = 16'b11111111_01100110;
		Dminus[398] = 16'b11111111_01100110;
		Dminus[399] = 16'b11111111_01100111;
		Dminus[400] = 16'b11111111_01100111;
		Dminus[401] = 16'b11111111_01101000;
		Dminus[402] = 16'b11111111_01101000;
		Dminus[403] = 16'b11111111_01101001;
		Dminus[404] = 16'b11111111_01101001;
		Dminus[405] = 16'b11111111_01101010;
		Dminus[406] = 16'b11111111_01101010;
		Dminus[407] = 16'b11111111_01101011;
		Dminus[408] = 16'b11111111_01101011;
		Dminus[409] = 16'b11111111_01101100;
		Dminus[410] = 16'b11111111_01101100;
		Dminus[411] = 16'b11111111_01101101;
		Dminus[412] = 16'b11111111_01101101;
		Dminus[413] = 16'b11111111_01101110;
		Dminus[414] = 16'b11111111_01101110;
		Dminus[415] = 16'b11111111_01101111;
		Dminus[416] = 16'b11111111_01101111;
		Dminus[417] = 16'b11111111_01110000;
		Dminus[418] = 16'b11111111_01110000;
		Dminus[419] = 16'b11111111_01110001;
		Dminus[420] = 16'b11111111_01110001;
		Dminus[421] = 16'b11111111_01110010;
		Dminus[422] = 16'b11111111_01110010;
		Dminus[423] = 16'b11111111_01110011;
		Dminus[424] = 16'b11111111_01110011;
		Dminus[425] = 16'b11111111_01110100;
		Dminus[426] = 16'b11111111_01110100;
		Dminus[427] = 16'b11111111_01110100;
		Dminus[428] = 16'b11111111_01110101;
		Dminus[429] = 16'b11111111_01110101;
		Dminus[430] = 16'b11111111_01110110;
		Dminus[431] = 16'b11111111_01110110;
		Dminus[432] = 16'b11111111_01110111;
		Dminus[433] = 16'b11111111_01110111;
		Dminus[434] = 16'b11111111_01111000;
		Dminus[435] = 16'b11111111_01111000;
		Dminus[436] = 16'b11111111_01111000;
		Dminus[437] = 16'b11111111_01111001;
		Dminus[438] = 16'b11111111_01111001;
		Dminus[439] = 16'b11111111_01111010;
		Dminus[440] = 16'b11111111_01111010;
		Dminus[441] = 16'b11111111_01111011;
		Dminus[442] = 16'b11111111_01111011;
		Dminus[443] = 16'b11111111_01111100;
		Dminus[444] = 16'b11111111_01111100;
		Dminus[445] = 16'b11111111_01111100;
		Dminus[446] = 16'b11111111_01111101;
		Dminus[447] = 16'b11111111_01111101;
		Dminus[448] = 16'b11111111_01111110;
		Dminus[449] = 16'b11111111_01111110;
		Dminus[450] = 16'b11111111_01111111;
		Dminus[451] = 16'b11111111_01111111;
		Dminus[452] = 16'b11111111_01111111;
		Dminus[453] = 16'b11111111_10000000;
		Dminus[454] = 16'b11111111_10000000;
		Dminus[455] = 16'b11111111_10000001;
		Dminus[456] = 16'b11111111_10000001;
		Dminus[457] = 16'b11111111_10000001;
		Dminus[458] = 16'b11111111_10000010;
		Dminus[459] = 16'b11111111_10000010;
		Dminus[460] = 16'b11111111_10000011;
		Dminus[461] = 16'b11111111_10000011;
		Dminus[462] = 16'b11111111_10000011;
		Dminus[463] = 16'b11111111_10000100;
		Dminus[464] = 16'b11111111_10000100;
		Dminus[465] = 16'b11111111_10000101;
		Dminus[466] = 16'b11111111_10000101;
		Dminus[467] = 16'b11111111_10000101;
		Dminus[468] = 16'b11111111_10000110;
		Dminus[469] = 16'b11111111_10000110;
		Dminus[470] = 16'b11111111_10000111;
		Dminus[471] = 16'b11111111_10000111;
		Dminus[472] = 16'b11111111_10000111;
		Dminus[473] = 16'b11111111_10001000;
		Dminus[474] = 16'b11111111_10001000;
		Dminus[475] = 16'b11111111_10001001;
		Dminus[476] = 16'b11111111_10001001;
		Dminus[477] = 16'b11111111_10001001;
		Dminus[478] = 16'b11111111_10001010;
		Dminus[479] = 16'b11111111_10001010;
		Dminus[480] = 16'b11111111_10001010;
		Dminus[481] = 16'b11111111_10001011;
		Dminus[482] = 16'b11111111_10001011;
		Dminus[483] = 16'b11111111_10001100;
		Dminus[484] = 16'b11111111_10001100;
		Dminus[485] = 16'b11111111_10001100;
		Dminus[486] = 16'b11111111_10001101;
		Dminus[487] = 16'b11111111_10001101;
		Dminus[488] = 16'b11111111_10001101;
		Dminus[489] = 16'b11111111_10001110;
		Dminus[490] = 16'b11111111_10001110;
		Dminus[491] = 16'b11111111_10001110;
		Dminus[492] = 16'b11111111_10001111;
		Dminus[493] = 16'b11111111_10001111;
		Dminus[494] = 16'b11111111_10010000;
		Dminus[495] = 16'b11111111_10010000;
		Dminus[496] = 16'b11111111_10010000;
		Dminus[497] = 16'b11111111_10010001;
		Dminus[498] = 16'b11111111_10010001;
		Dminus[499] = 16'b11111111_10010001;
		Dminus[500] = 16'b11111111_10010010;
		Dminus[501] = 16'b11111111_10010010;
		Dminus[502] = 16'b11111111_10010010;
		Dminus[503] = 16'b11111111_10010011;
		Dminus[504] = 16'b11111111_10010011;
		Dminus[505] = 16'b11111111_10010011;
		Dminus[506] = 16'b11111111_10010100;
		Dminus[507] = 16'b11111111_10010100;
		Dminus[508] = 16'b11111111_10010100;
		Dminus[509] = 16'b11111111_10010101;
		Dminus[510] = 16'b11111111_10010101;
		Dminus[511] = 16'b11111111_10010101;
		Dplus[1] = 16'b00000001_00000000;
		Dplus[2] = 16'b00000000_11111111;
		Dplus[3] = 16'b00000000_11111111;
		Dplus[4] = 16'b00000000_11111110;
		Dplus[5] = 16'b00000000_11111110;
		Dplus[6] = 16'b00000000_11111101;
		Dplus[7] = 16'b00000000_11111101;
		Dplus[8] = 16'b00000000_11111100;
		Dplus[9] = 16'b00000000_11111100;
		Dplus[10] = 16'b00000000_11111011;
		Dplus[11] = 16'b00000000_11111011;
		Dplus[12] = 16'b00000000_11111010;
		Dplus[13] = 16'b00000000_11111010;
		Dplus[14] = 16'b00000000_11111001;
		Dplus[15] = 16'b00000000_11111001;
		Dplus[16] = 16'b00000000_11111000;
		Dplus[17] = 16'b00000000_11111000;
		Dplus[18] = 16'b00000000_11110111;
		Dplus[19] = 16'b00000000_11110111;
		Dplus[20] = 16'b00000000_11110110;
		Dplus[21] = 16'b00000000_11110110;
		Dplus[22] = 16'b00000000_11110101;
		Dplus[23] = 16'b00000000_11110101;
		Dplus[24] = 16'b00000000_11110100;
		Dplus[25] = 16'b00000000_11110100;
		Dplus[26] = 16'b00000000_11110011;
		Dplus[27] = 16'b00000000_11110011;
		Dplus[28] = 16'b00000000_11110010;
		Dplus[29] = 16'b00000000_11110010;
		Dplus[30] = 16'b00000000_11110001;
		Dplus[31] = 16'b00000000_11110001;
		Dplus[32] = 16'b00000000_11110000;
		Dplus[33] = 16'b00000000_11110000;
		Dplus[34] = 16'b00000000_11101111;
		Dplus[35] = 16'b00000000_11101111;
		Dplus[36] = 16'b00000000_11101110;
		Dplus[37] = 16'b00000000_11101110;
		Dplus[38] = 16'b00000000_11101101;
		Dplus[39] = 16'b00000000_11101101;
		Dplus[40] = 16'b00000000_11101101;
		Dplus[41] = 16'b00000000_11101100;
		Dplus[42] = 16'b00000000_11101100;
		Dplus[43] = 16'b00000000_11101011;
		Dplus[44] = 16'b00000000_11101011;
		Dplus[45] = 16'b00000000_11101010;
		Dplus[46] = 16'b00000000_11101010;
		Dplus[47] = 16'b00000000_11101001;
		Dplus[48] = 16'b00000000_11101001;
		Dplus[49] = 16'b00000000_11101000;
		Dplus[50] = 16'b00000000_11101000;
		Dplus[51] = 16'b00000000_11100111;
		Dplus[52] = 16'b00000000_11100111;
		Dplus[53] = 16'b00000000_11100110;
		Dplus[54] = 16'b00000000_11100110;
		Dplus[55] = 16'b00000000_11100110;
		Dplus[56] = 16'b00000000_11100101;
		Dplus[57] = 16'b00000000_11100101;
		Dplus[58] = 16'b00000000_11100100;
		Dplus[59] = 16'b00000000_11100100;
		Dplus[60] = 16'b00000000_11100011;
		Dplus[61] = 16'b00000000_11100011;
		Dplus[62] = 16'b00000000_11100010;
		Dplus[63] = 16'b00000000_11100010;
		Dplus[64] = 16'b00000000_11100001;
		Dplus[65] = 16'b00000000_11100001;
		Dplus[66] = 16'b00000000_11100000;
		Dplus[67] = 16'b00000000_11100000;
		Dplus[68] = 16'b00000000_11100000;
		Dplus[69] = 16'b00000000_11011111;
		Dplus[70] = 16'b00000000_11011111;
		Dplus[71] = 16'b00000000_11011110;
		Dplus[72] = 16'b00000000_11011110;
		Dplus[73] = 16'b00000000_11011101;
		Dplus[74] = 16'b00000000_11011101;
		Dplus[75] = 16'b00000000_11011100;
		Dplus[76] = 16'b00000000_11011100;
		Dplus[77] = 16'b00000000_11011100;
		Dplus[78] = 16'b00000000_11011011;
		Dplus[79] = 16'b00000000_11011011;
		Dplus[80] = 16'b00000000_11011010;
		Dplus[81] = 16'b00000000_11011010;
		Dplus[82] = 16'b00000000_11011001;
		Dplus[83] = 16'b00000000_11011001;
		Dplus[84] = 16'b00000000_11011000;
		Dplus[85] = 16'b00000000_11011000;
		Dplus[86] = 16'b00000000_11010111;
		Dplus[87] = 16'b00000000_11010111;
		Dplus[88] = 16'b00000000_11010111;
		Dplus[89] = 16'b00000000_11010110;
		Dplus[90] = 16'b00000000_11010110;
		Dplus[91] = 16'b00000000_11010101;
		Dplus[92] = 16'b00000000_11010101;
		Dplus[93] = 16'b00000000_11010100;
		Dplus[94] = 16'b00000000_11010100;
		Dplus[95] = 16'b00000000_11010100;
		Dplus[96] = 16'b00000000_11010011;
		Dplus[97] = 16'b00000000_11010011;
		Dplus[98] = 16'b00000000_11010010;
		Dplus[99] = 16'b00000000_11010010;
		Dplus[100] = 16'b00000000_11010001;
		Dplus[101] = 16'b00000000_11010001;
		Dplus[102] = 16'b00000000_11010001;
		Dplus[103] = 16'b00000000_11010000;
		Dplus[104] = 16'b00000000_11010000;
		Dplus[105] = 16'b00000000_11001111;
		Dplus[106] = 16'b00000000_11001111;
		Dplus[107] = 16'b00000000_11001110;
		Dplus[108] = 16'b00000000_11001110;
		Dplus[109] = 16'b00000000_11001110;
		Dplus[110] = 16'b00000000_11001101;
		Dplus[111] = 16'b00000000_11001101;
		Dplus[112] = 16'b00000000_11001100;
		Dplus[113] = 16'b00000000_11001100;
		Dplus[114] = 16'b00000000_11001011;
		Dplus[115] = 16'b00000000_11001011;
		Dplus[116] = 16'b00000000_11001011;
		Dplus[117] = 16'b00000000_11001010;
		Dplus[118] = 16'b00000000_11001010;
		Dplus[119] = 16'b00000000_11001001;
		Dplus[120] = 16'b00000000_11001001;
		Dplus[121] = 16'b00000000_11001000;
		Dplus[122] = 16'b00000000_11001000;
		Dplus[123] = 16'b00000000_11001000;
		Dplus[124] = 16'b00000000_11000111;
		Dplus[125] = 16'b00000000_11000111;
		Dplus[126] = 16'b00000000_11000110;
		Dplus[127] = 16'b00000000_11000110;
		Dplus[128] = 16'b00000000_11000110;
		Dplus[129] = 16'b00000000_11000101;
		Dplus[130] = 16'b00000000_11000101;
		Dplus[131] = 16'b00000000_11000100;
		Dplus[132] = 16'b00000000_11000100;
		Dplus[133] = 16'b00000000_11000011;
		Dplus[134] = 16'b00000000_11000011;
		Dplus[135] = 16'b00000000_11000011;
		Dplus[136] = 16'b00000000_11000010;
		Dplus[137] = 16'b00000000_11000010;
		Dplus[138] = 16'b00000000_11000001;
		Dplus[139] = 16'b00000000_11000001;
		Dplus[140] = 16'b00000000_11000001;
		Dplus[141] = 16'b00000000_11000000;
		Dplus[142] = 16'b00000000_11000000;
		Dplus[143] = 16'b00000000_10111111;
		Dplus[144] = 16'b00000000_10111111;
		Dplus[145] = 16'b00000000_10111111;
		Dplus[146] = 16'b00000000_10111110;
		Dplus[147] = 16'b00000000_10111110;
		Dplus[148] = 16'b00000000_10111101;
		Dplus[149] = 16'b00000000_10111101;
		Dplus[150] = 16'b00000000_10111101;
		Dplus[151] = 16'b00000000_10111100;
		Dplus[152] = 16'b00000000_10111100;
		Dplus[153] = 16'b00000000_10111011;
		Dplus[154] = 16'b00000000_10111011;
		Dplus[155] = 16'b00000000_10111011;
		Dplus[156] = 16'b00000000_10111010;
		Dplus[157] = 16'b00000000_10111010;
		Dplus[158] = 16'b00000000_10111001;
		Dplus[159] = 16'b00000000_10111001;
		Dplus[160] = 16'b00000000_10111001;
		Dplus[161] = 16'b00000000_10111000;
		Dplus[162] = 16'b00000000_10111000;
		Dplus[163] = 16'b00000000_10110111;
		Dplus[164] = 16'b00000000_10110111;
		Dplus[165] = 16'b00000000_10110111;
		Dplus[166] = 16'b00000000_10110110;
		Dplus[167] = 16'b00000000_10110110;
		Dplus[168] = 16'b00000000_10110101;
		Dplus[169] = 16'b00000000_10110101;
		Dplus[170] = 16'b00000000_10110101;
		Dplus[171] = 16'b00000000_10110100;
		Dplus[172] = 16'b00000000_10110100;
		Dplus[173] = 16'b00000000_10110100;
		Dplus[174] = 16'b00000000_10110011;
		Dplus[175] = 16'b00000000_10110011;
		Dplus[176] = 16'b00000000_10110010;
		Dplus[177] = 16'b00000000_10110010;
		Dplus[178] = 16'b00000000_10110010;
		Dplus[179] = 16'b00000000_10110001;
		Dplus[180] = 16'b00000000_10110001;
		Dplus[181] = 16'b00000000_10110000;
		Dplus[182] = 16'b00000000_10110000;
		Dplus[183] = 16'b00000000_10110000;
		Dplus[184] = 16'b00000000_10101111;
		Dplus[185] = 16'b00000000_10101111;
		Dplus[186] = 16'b00000000_10101111;
		Dplus[187] = 16'b00000000_10101110;
		Dplus[188] = 16'b00000000_10101110;
		Dplus[189] = 16'b00000000_10101101;
		Dplus[190] = 16'b00000000_10101101;
		Dplus[191] = 16'b00000000_10101101;
		Dplus[192] = 16'b00000000_10101100;
		Dplus[193] = 16'b00000000_10101100;
		Dplus[194] = 16'b00000000_10101100;
		Dplus[195] = 16'b00000000_10101011;
		Dplus[196] = 16'b00000000_10101011;
		Dplus[197] = 16'b00000000_10101010;
		Dplus[198] = 16'b00000000_10101010;
		Dplus[199] = 16'b00000000_10101010;
		Dplus[200] = 16'b00000000_10101001;
		Dplus[201] = 16'b00000000_10101001;
		Dplus[202] = 16'b00000000_10101001;
		Dplus[203] = 16'b00000000_10101000;
		Dplus[204] = 16'b00000000_10101000;
		Dplus[205] = 16'b00000000_10101000;
		Dplus[206] = 16'b00000000_10100111;
		Dplus[207] = 16'b00000000_10100111;
		Dplus[208] = 16'b00000000_10100110;
		Dplus[209] = 16'b00000000_10100110;
		Dplus[210] = 16'b00000000_10100110;
		Dplus[211] = 16'b00000000_10100101;
		Dplus[212] = 16'b00000000_10100101;
		Dplus[213] = 16'b00000000_10100101;
		Dplus[214] = 16'b00000000_10100100;
		Dplus[215] = 16'b00000000_10100100;
		Dplus[216] = 16'b00000000_10100100;
		Dplus[217] = 16'b00000000_10100011;
		Dplus[218] = 16'b00000000_10100011;
		Dplus[219] = 16'b00000000_10100011;
		Dplus[220] = 16'b00000000_10100010;
		Dplus[221] = 16'b00000000_10100010;
		Dplus[222] = 16'b00000000_10100001;
		Dplus[223] = 16'b00000000_10100001;
		Dplus[224] = 16'b00000000_10100001;
		Dplus[225] = 16'b00000000_10100000;
		Dplus[226] = 16'b00000000_10100000;
		Dplus[227] = 16'b00000000_10100000;
		Dplus[228] = 16'b00000000_10011111;
		Dplus[229] = 16'b00000000_10011111;
		Dplus[230] = 16'b00000000_10011111;
		Dplus[231] = 16'b00000000_10011110;
		Dplus[232] = 16'b00000000_10011110;
		Dplus[233] = 16'b00000000_10011110;
		Dplus[234] = 16'b00000000_10011101;
		Dplus[235] = 16'b00000000_10011101;
		Dplus[236] = 16'b00000000_10011101;
		Dplus[237] = 16'b00000000_10011100;
		Dplus[238] = 16'b00000000_10011100;
		Dplus[239] = 16'b00000000_10011100;
		Dplus[240] = 16'b00000000_10011011;
		Dplus[241] = 16'b00000000_10011011;
		Dplus[242] = 16'b00000000_10011010;
		Dplus[243] = 16'b00000000_10011010;
		Dplus[244] = 16'b00000000_10011010;
		Dplus[245] = 16'b00000000_10011001;
		Dplus[246] = 16'b00000000_10011001;
		Dplus[247] = 16'b00000000_10011001;
		Dplus[248] = 16'b00000000_10011000;
		Dplus[249] = 16'b00000000_10011000;
		Dplus[250] = 16'b00000000_10011000;
		Dplus[251] = 16'b00000000_10010111;
		Dplus[252] = 16'b00000000_10010111;
		Dplus[253] = 16'b00000000_10010111;
		Dplus[254] = 16'b00000000_10010110;
		Dplus[255] = 16'b00000000_10010110;
		Dplus[256] = 16'b00000000_10010110;
		Dplus[257] = 16'b00000000_10010101;
		Dplus[258] = 16'b00000000_10010101;
		Dplus[259] = 16'b00000000_10010101;
		Dplus[260] = 16'b00000000_10010100;
		Dplus[261] = 16'b00000000_10010100;
		Dplus[262] = 16'b00000000_10010100;
		Dplus[263] = 16'b00000000_10010011;
		Dplus[264] = 16'b00000000_10010011;
		Dplus[265] = 16'b00000000_10010011;
		Dplus[266] = 16'b00000000_10010010;
		Dplus[267] = 16'b00000000_10010010;
		Dplus[268] = 16'b00000000_10010010;
		Dplus[269] = 16'b00000000_10010001;
		Dplus[270] = 16'b00000000_10010001;
		Dplus[271] = 16'b00000000_10010001;
		Dplus[272] = 16'b00000000_10010000;
		Dplus[273] = 16'b00000000_10010000;
		Dplus[274] = 16'b00000000_10010000;
		Dplus[275] = 16'b00000000_10010000;
		Dplus[276] = 16'b00000000_10001111;
		Dplus[277] = 16'b00000000_10001111;
		Dplus[278] = 16'b00000000_10001111;
		Dplus[279] = 16'b00000000_10001110;
		Dplus[280] = 16'b00000000_10001110;
		Dplus[281] = 16'b00000000_10001110;
		Dplus[282] = 16'b00000000_10001101;
		Dplus[283] = 16'b00000000_10001101;
		Dplus[284] = 16'b00000000_10001101;
		Dplus[285] = 16'b00000000_10001100;
		Dplus[286] = 16'b00000000_10001100;
		Dplus[287] = 16'b00000000_10001100;
		Dplus[288] = 16'b00000000_10001011;
		Dplus[289] = 16'b00000000_10001011;
		Dplus[290] = 16'b00000000_10001011;
		Dplus[291] = 16'b00000000_10001010;
		Dplus[292] = 16'b00000000_10001010;
		Dplus[293] = 16'b00000000_10001010;
		Dplus[294] = 16'b00000000_10001010;
		Dplus[295] = 16'b00000000_10001001;
		Dplus[296] = 16'b00000000_10001001;
		Dplus[297] = 16'b00000000_10001001;
		Dplus[298] = 16'b00000000_10001000;
		Dplus[299] = 16'b00000000_10001000;
		Dplus[300] = 16'b00000000_10001000;
		Dplus[301] = 16'b00000000_10000111;
		Dplus[302] = 16'b00000000_10000111;
		Dplus[303] = 16'b00000000_10000111;
		Dplus[304] = 16'b00000000_10000110;
		Dplus[305] = 16'b00000000_10000110;
		Dplus[306] = 16'b00000000_10000110;
		Dplus[307] = 16'b00000000_10000110;
		Dplus[308] = 16'b00000000_10000101;
		Dplus[309] = 16'b00000000_10000101;
		Dplus[310] = 16'b00000000_10000101;
		Dplus[311] = 16'b00000000_10000100;
		Dplus[312] = 16'b00000000_10000100;
		Dplus[313] = 16'b00000000_10000100;
		Dplus[314] = 16'b00000000_10000011;
		Dplus[315] = 16'b00000000_10000011;
		Dplus[316] = 16'b00000000_10000011;
		Dplus[317] = 16'b00000000_10000011;
		Dplus[318] = 16'b00000000_10000010;
		Dplus[319] = 16'b00000000_10000010;
		Dplus[320] = 16'b00000000_10000010;
		Dplus[321] = 16'b00000000_10000001;
		Dplus[322] = 16'b00000000_10000001;
		Dplus[323] = 16'b00000000_10000001;
		Dplus[324] = 16'b00000000_10000000;
		Dplus[325] = 16'b00000000_10000000;
		Dplus[326] = 16'b00000000_10000000;
		Dplus[327] = 16'b00000000_10000000;
		Dplus[328] = 16'b00000000_01111111;
		Dplus[329] = 16'b00000000_01111111;
		Dplus[330] = 16'b00000000_01111111;
		Dplus[331] = 16'b00000000_01111110;
		Dplus[332] = 16'b00000000_01111110;
		Dplus[333] = 16'b00000000_01111110;
		Dplus[334] = 16'b00000000_01111110;
		Dplus[335] = 16'b00000000_01111101;
		Dplus[336] = 16'b00000000_01111101;
		Dplus[337] = 16'b00000000_01111101;
		Dplus[338] = 16'b00000000_01111100;
		Dplus[339] = 16'b00000000_01111100;
		Dplus[340] = 16'b00000000_01111100;
		Dplus[341] = 16'b00000000_01111100;
		Dplus[342] = 16'b00000000_01111011;
		Dplus[343] = 16'b00000000_01111011;
		Dplus[344] = 16'b00000000_01111011;
		Dplus[345] = 16'b00000000_01111010;
		Dplus[346] = 16'b00000000_01111010;
		Dplus[347] = 16'b00000000_01111010;
		Dplus[348] = 16'b00000000_01111010;
		Dplus[349] = 16'b00000000_01111001;
		Dplus[350] = 16'b00000000_01111001;
		Dplus[351] = 16'b00000000_01111001;
		Dplus[352] = 16'b00000000_01111000;
		Dplus[353] = 16'b00000000_01111000;
		Dplus[354] = 16'b00000000_01111000;
		Dplus[355] = 16'b00000000_01111000;
		Dplus[356] = 16'b00000000_01110111;
		Dplus[357] = 16'b00000000_01110111;
		Dplus[358] = 16'b00000000_01110111;
		Dplus[359] = 16'b00000000_01110111;
		Dplus[360] = 16'b00000000_01110110;
		Dplus[361] = 16'b00000000_01110110;
		Dplus[362] = 16'b00000000_01110110;
		Dplus[363] = 16'b00000000_01110101;
		Dplus[364] = 16'b00000000_01110101;
		Dplus[365] = 16'b00000000_01110101;
		Dplus[366] = 16'b00000000_01110101;
		Dplus[367] = 16'b00000000_01110100;
		Dplus[368] = 16'b00000000_01110100;
		Dplus[369] = 16'b00000000_01110100;
		Dplus[370] = 16'b00000000_01110100;
		Dplus[371] = 16'b00000000_01110011;
		Dplus[372] = 16'b00000000_01110011;
		Dplus[373] = 16'b00000000_01110011;
		Dplus[374] = 16'b00000000_01110010;
		Dplus[375] = 16'b00000000_01110010;
		Dplus[376] = 16'b00000000_01110010;
		Dplus[377] = 16'b00000000_01110010;
		Dplus[378] = 16'b00000000_01110001;
		Dplus[379] = 16'b00000000_01110001;
		Dplus[380] = 16'b00000000_01110001;
		Dplus[381] = 16'b00000000_01110001;
		Dplus[382] = 16'b00000000_01110000;
		Dplus[383] = 16'b00000000_01110000;
		Dplus[384] = 16'b00000000_01110000;
		Dplus[385] = 16'b00000000_01110000;
		Dplus[386] = 16'b00000000_01101111;
		Dplus[387] = 16'b00000000_01101111;
		Dplus[388] = 16'b00000000_01101111;
		Dplus[389] = 16'b00000000_01101111;
		Dplus[390] = 16'b00000000_01101110;
		Dplus[391] = 16'b00000000_01101110;
		Dplus[392] = 16'b00000000_01101110;
		Dplus[393] = 16'b00000000_01101101;
		Dplus[394] = 16'b00000000_01101101;
		Dplus[395] = 16'b00000000_01101101;
		Dplus[396] = 16'b00000000_01101101;
		Dplus[397] = 16'b00000000_01101100;
		Dplus[398] = 16'b00000000_01101100;
		Dplus[399] = 16'b00000000_01101100;
		Dplus[400] = 16'b00000000_01101100;
		Dplus[401] = 16'b00000000_01101011;
		Dplus[402] = 16'b00000000_01101011;
		Dplus[403] = 16'b00000000_01101011;
		Dplus[404] = 16'b00000000_01101011;
		Dplus[405] = 16'b00000000_01101010;
		Dplus[406] = 16'b00000000_01101010;
		Dplus[407] = 16'b00000000_01101010;
		Dplus[408] = 16'b00000000_01101010;
		Dplus[409] = 16'b00000000_01101001;
		Dplus[410] = 16'b00000000_01101001;
		Dplus[411] = 16'b00000000_01101001;
		Dplus[412] = 16'b00000000_01101001;
		Dplus[413] = 16'b00000000_01101000;
		Dplus[414] = 16'b00000000_01101000;
		Dplus[415] = 16'b00000000_01101000;
		Dplus[416] = 16'b00000000_01101000;
		Dplus[417] = 16'b00000000_01100111;
		Dplus[418] = 16'b00000000_01100111;
		Dplus[419] = 16'b00000000_01100111;
		Dplus[420] = 16'b00000000_01100111;
		Dplus[421] = 16'b00000000_01100110;
		Dplus[422] = 16'b00000000_01100110;
		Dplus[423] = 16'b00000000_01100110;
		Dplus[424] = 16'b00000000_01100110;
		Dplus[425] = 16'b00000000_01100110;
		Dplus[426] = 16'b00000000_01100101;
		Dplus[427] = 16'b00000000_01100101;
		Dplus[428] = 16'b00000000_01100101;
		Dplus[429] = 16'b00000000_01100101;
		Dplus[430] = 16'b00000000_01100100;
		Dplus[431] = 16'b00000000_01100100;
		Dplus[432] = 16'b00000000_01100100;
		Dplus[433] = 16'b00000000_01100100;
		Dplus[434] = 16'b00000000_01100011;
		Dplus[435] = 16'b00000000_01100011;
		Dplus[436] = 16'b00000000_01100011;
		Dplus[437] = 16'b00000000_01100011;
		Dplus[438] = 16'b00000000_01100010;
		Dplus[439] = 16'b00000000_01100010;
		Dplus[440] = 16'b00000000_01100010;
		Dplus[441] = 16'b00000000_01100010;
		Dplus[442] = 16'b00000000_01100010;
		Dplus[443] = 16'b00000000_01100001;
		Dplus[444] = 16'b00000000_01100001;
		Dplus[445] = 16'b00000000_01100001;
		Dplus[446] = 16'b00000000_01100001;
		Dplus[447] = 16'b00000000_01100000;
		Dplus[448] = 16'b00000000_01100000;
		Dplus[449] = 16'b00000000_01100000;
		Dplus[450] = 16'b00000000_01100000;
		Dplus[451] = 16'b00000000_01011111;
		Dplus[452] = 16'b00000000_01011111;
		Dplus[453] = 16'b00000000_01011111;
		Dplus[454] = 16'b00000000_01011111;
		Dplus[455] = 16'b00000000_01011111;
		Dplus[456] = 16'b00000000_01011110;
		Dplus[457] = 16'b00000000_01011110;
		Dplus[458] = 16'b00000000_01011110;
		Dplus[459] = 16'b00000000_01011110;
		Dplus[460] = 16'b00000000_01011101;
		Dplus[461] = 16'b00000000_01011101;
		Dplus[462] = 16'b00000000_01011101;
		Dplus[463] = 16'b00000000_01011101;
		Dplus[464] = 16'b00000000_01011101;
		Dplus[465] = 16'b00000000_01011100;
		Dplus[466] = 16'b00000000_01011100;
		Dplus[467] = 16'b00000000_01011100;
		Dplus[468] = 16'b00000000_01011100;
		Dplus[469] = 16'b00000000_01011011;
		Dplus[470] = 16'b00000000_01011011;
		Dplus[471] = 16'b00000000_01011011;
		Dplus[472] = 16'b00000000_01011011;
		Dplus[473] = 16'b00000000_01011011;
		Dplus[474] = 16'b00000000_01011010;
		Dplus[475] = 16'b00000000_01011010;
		Dplus[476] = 16'b00000000_01011010;
		Dplus[477] = 16'b00000000_01011010;
		Dplus[478] = 16'b00000000_01011001;
		Dplus[479] = 16'b00000000_01011001;
		Dplus[480] = 16'b00000000_01011001;
		Dplus[481] = 16'b00000000_01011001;
		Dplus[482] = 16'b00000000_01011001;
		Dplus[483] = 16'b00000000_01011000;
		Dplus[484] = 16'b00000000_01011000;
		Dplus[485] = 16'b00000000_01011000;
		Dplus[486] = 16'b00000000_01011000;
		Dplus[487] = 16'b00000000_01011000;
		Dplus[488] = 16'b00000000_01010111;
		Dplus[489] = 16'b00000000_01010111;
		Dplus[490] = 16'b00000000_01010111;
		Dplus[491] = 16'b00000000_01010111;
		Dplus[492] = 16'b00000000_01010111;
		Dplus[493] = 16'b00000000_01010110;
		Dplus[494] = 16'b00000000_01010110;
		Dplus[495] = 16'b00000000_01010110;
		Dplus[496] = 16'b00000000_01010110;
		Dplus[497] = 16'b00000000_01010101;
		Dplus[498] = 16'b00000000_01010101;
		Dplus[499] = 16'b00000000_01010101;
		Dplus[500] = 16'b00000000_01010101;
		Dplus[501] = 16'b00000000_01010101;
		Dplus[502] = 16'b00000000_01010100;
		Dplus[503] = 16'b00000000_01010100;
		Dplus[504] = 16'b00000000_01010100;
		Dplus[505] = 16'b00000000_01010100;
		Dplus[506] = 16'b00000000_01010100;
		Dplus[507] = 16'b00000000_01010011;
		Dplus[508] = 16'b00000000_01010011;
		Dplus[509] = 16'b00000000_01010011;
		Dplus[510] = 16'b00000000_01010011;
		Dplus[511] = 16'b00000000_01010011;
		DplusInteger[2] = 16'b00000000_01010010;
		DplusInteger[3] = 16'b00000000_00101100;
		DplusInteger[4] = 16'b00000000_00010110;
		DplusInteger[5] = 16'b00000000_00001011;
		DplusInteger[6] = 16'b00000000_00000110;
		DplusInteger[7] = 16'b00000000_00000011;
		DplusInteger[8] = 16'b00000000_00000001;
		DplusInteger[9] = 16'b00000000_00000001;
		DplusInteger[10] = 16'b00000000_00000000;
		DplusInteger[11] = 16'b00000000_00000000;
		DplusInteger[12] = 16'b00000000_00000000;
		DplusInteger[13] = 16'b00000000_00000000;
		DplusInteger[14] = 16'b00000000_00000000;
		DplusInteger[15] = 16'b00000000_00000000;
		DplusInteger[16] = 16'b00000000_00000000;
		DplusInteger[17] = 16'b00000000_00000000;
		DplusInteger[18] = 16'b00000000_00000000;
		DplusInteger[19] = 16'b00000000_00000000;
		DplusInteger[20] = 16'b00000000_00000000;
		DplusInteger[21] = 16'b00000000_00000000;
		DplusInteger[22] = 16'b00000000_00000000;
		DplusInteger[23] = 16'b00000000_00000000;
		DplusInteger[24] = 16'b00000000_00000000;
		DplusInteger[25] = 16'b00000000_00000000;
		DplusInteger[26] = 16'b00000000_00000000;
		DplusInteger[27] = 16'b00000000_00000000;
		DplusInteger[28] = 16'b00000000_00000000;
		DplusInteger[29] = 16'b00000000_00000000;
		DplusInteger[30] = 16'b00000000_00000000;
		DplusInteger[31] = 16'b00000000_00000000;
		DplusInteger[32] = 16'b00000000_00000000;
		DplusInteger[33] = 16'b00000000_00000000;
		DplusInteger[34] = 16'b00000000_00000000;
		DplusInteger[35] = 16'b00000000_00000000;
		DplusInteger[36] = 16'b00000000_00000000;
		DplusInteger[37] = 16'b00000000_00000000;
		DplusInteger[38] = 16'b00000000_00000000;
		DplusInteger[39] = 16'b00000000_00000000;
		DplusInteger[40] = 16'b00000000_00000000;
		DplusInteger[41] = 16'b00000000_00000000;
		DplusInteger[42] = 16'b00000000_00000000;
		DplusInteger[43] = 16'b00000000_00000000;
		DplusInteger[44] = 16'b00000000_00000000;
		DplusInteger[45] = 16'b00000000_00000000;
		DplusInteger[46] = 16'b00000000_00000000;
		DplusInteger[47] = 16'b00000000_00000000;
		DplusInteger[48] = 16'b00000000_00000000;
		DplusInteger[49] = 16'b00000000_00000000;
		DplusInteger[50] = 16'b00000000_00000000;
		DplusInteger[51] = 16'b00000000_00000000;
		DplusInteger[52] = 16'b00000000_00000000;
		DplusInteger[53] = 16'b00000000_00000000;
		DplusInteger[54] = 16'b00000000_00000000;
		DplusInteger[55] = 16'b00000000_00000000;
		DplusInteger[56] = 16'b00000000_00000000;
		DplusInteger[57] = 16'b00000000_00000000;
		DplusInteger[58] = 16'b00000000_00000000;
		DplusInteger[59] = 16'b00000000_00000000;
		DplusInteger[60] = 16'b00000000_00000000;
		DplusInteger[61] = 16'b00000000_00000000;
		DplusInteger[62] = 16'b00000000_00000000;
		DplusInteger[63] = 16'b00000000_00000000;
		DplusInteger[64] = 16'b00000000_00000000;
		DplusInteger[65] = 16'b00000000_00000000;
		DplusInteger[66] = 16'b00000000_00000000;
		DplusInteger[67] = 16'b00000000_00000000;
		DplusInteger[68] = 16'b00000000_00000000;
		DplusInteger[69] = 16'b00000000_00000000;
		DplusInteger[70] = 16'b00000000_00000000;
		DplusInteger[71] = 16'b00000000_00000000;
		DplusInteger[72] = 16'b00000000_00000000;
		DplusInteger[73] = 16'b00000000_00000000;
		DplusInteger[74] = 16'b00000000_00000000;
		DplusInteger[75] = 16'b00000000_00000000;
		DplusInteger[76] = 16'b00000000_00000000;
		DplusInteger[77] = 16'b00000000_00000000;
		DplusInteger[78] = 16'b00000000_00000000;
		DplusInteger[79] = 16'b00000000_00000000;
		DplusInteger[80] = 16'b00000000_00000000;
		DplusInteger[81] = 16'b00000000_00000000;
		DplusInteger[82] = 16'b00000000_00000000;
		DplusInteger[83] = 16'b00000000_00000000;
		DplusInteger[84] = 16'b00000000_00000000;
		DplusInteger[85] = 16'b00000000_00000000;
		DplusInteger[86] = 16'b00000000_00000000;
		DplusInteger[87] = 16'b00000000_00000000;
		DplusInteger[88] = 16'b00000000_00000000;
		DplusInteger[89] = 16'b00000000_00000000;
		DplusInteger[90] = 16'b00000000_00000000;
		DplusInteger[91] = 16'b00000000_00000000;
		DplusInteger[92] = 16'b00000000_00000000;
		DplusInteger[93] = 16'b00000000_00000000;
		DplusInteger[94] = 16'b00000000_00000000;
		DplusInteger[95] = 16'b00000000_00000000;
		DplusInteger[96] = 16'b00000000_00000000;
		DplusInteger[97] = 16'b00000000_00000000;
		DplusInteger[98] = 16'b00000000_00000000;
		DplusInteger[99] = 16'b00000000_00000000;
		DplusInteger[100] = 16'b00000000_00000000;
		DplusInteger[101] = 16'b00000000_00000000;
		DplusInteger[102] = 16'b00000000_00000000;
		DplusInteger[103] = 16'b00000000_00000000;
		DplusInteger[104] = 16'b00000000_00000000;
		DplusInteger[105] = 16'b00000000_00000000;
		DplusInteger[106] = 16'b00000000_00000000;
		DplusInteger[107] = 16'b00000000_00000000;
		DplusInteger[108] = 16'b00000000_00000000;
		DplusInteger[109] = 16'b00000000_00000000;
		DplusInteger[110] = 16'b00000000_00000000;
		DplusInteger[111] = 16'b00000000_00000000;
		DplusInteger[112] = 16'b00000000_00000000;
		DplusInteger[113] = 16'b00000000_00000000;
		DplusInteger[114] = 16'b00000000_00000000;
		DplusInteger[115] = 16'b00000000_00000000;
		DplusInteger[116] = 16'b00000000_00000000;
		DplusInteger[117] = 16'b00000000_00000000;
		DplusInteger[118] = 16'b00000000_00000000;
		DplusInteger[119] = 16'b00000000_00000000;
		DplusInteger[120] = 16'b00000000_00000000;
		DplusInteger[121] = 16'b00000000_00000000;
		DplusInteger[122] = 16'b00000000_00000000;
		DplusInteger[123] = 16'b00000000_00000000;
		DplusInteger[124] = 16'b00000000_00000000;
		DplusInteger[125] = 16'b00000000_00000000;
		DplusInteger[126] = 16'b00000000_00000000;
		DplusInteger[127] = 16'b00000000_00000000;
		DminusInteger[2] = 16'b11111111_10010110;
		DminusInteger[3] = 16'b11111111_11001111;
		DminusInteger[4] = 16'b11111111_11101000;
		DminusInteger[5] = 16'b11111111_11110100;
		DminusInteger[6] = 16'b11111111_11111010;
		DminusInteger[7] = 16'b11111111_11111101;
		DminusInteger[8] = 16'b11111111_11111111;
		DminusInteger[9] = 16'b11111111_11111111;
		DminusInteger[10] = 16'b00000000_00000000;
		DminusInteger[11] = 16'b00000000_00000000;
		DminusInteger[12] = 16'b00000000_00000000;
		DminusInteger[13] = 16'b00000000_00000000;
		DminusInteger[14] = 16'b00000000_00000000;
		DminusInteger[15] = 16'b00000000_00000000;
		DminusInteger[16] = 16'b00000000_00000000;
		DminusInteger[17] = 16'b00000000_00000000;
		DminusInteger[18] = 16'b00000000_00000000;
		DminusInteger[19] = 16'b00000000_00000000;
		DminusInteger[20] = 16'b00000000_00000000;
		DminusInteger[21] = 16'b00000000_00000000;
		DminusInteger[22] = 16'b00000000_00000000;
		DminusInteger[23] = 16'b00000000_00000000;
		DminusInteger[24] = 16'b00000000_00000000;
		DminusInteger[25] = 16'b00000000_00000000;
		DminusInteger[26] = 16'b00000000_00000000;
		DminusInteger[27] = 16'b00000000_00000000;
		DminusInteger[28] = 16'b00000000_00000000;
		DminusInteger[29] = 16'b00000000_00000000;
		DminusInteger[30] = 16'b00000000_00000000;
		DminusInteger[31] = 16'b00000000_00000000;
		DminusInteger[32] = 16'b00000000_00000000;
		DminusInteger[33] = 16'b00000000_00000000;
		DminusInteger[34] = 16'b00000000_00000000;
		DminusInteger[35] = 16'b00000000_00000000;
		DminusInteger[36] = 16'b00000000_00000000;
		DminusInteger[37] = 16'b00000000_00000000;
		DminusInteger[38] = 16'b00000000_00000000;
		DminusInteger[39] = 16'b00000000_00000000;
		DminusInteger[40] = 16'b00000000_00000000;
		DminusInteger[41] = 16'b00000000_00000000;
		DminusInteger[42] = 16'b00000000_00000000;
		DminusInteger[43] = 16'b00000000_00000000;
		DminusInteger[44] = 16'b00000000_00000000;
		DminusInteger[45] = 16'b00000000_00000000;
		DminusInteger[46] = 16'b00000000_00000000;
		DminusInteger[47] = 16'b00000000_00000000;
		DminusInteger[48] = 16'b00000000_00000000;
		DminusInteger[49] = 16'b00000000_00000000;
		DminusInteger[50] = 16'b00000000_00000000;
		DminusInteger[51] = 16'b00000000_00000000;
		DminusInteger[52] = 16'b00000000_00000000;
		DminusInteger[53] = 16'b00000000_00000000;
		DminusInteger[54] = 16'b00000000_00000000;
		DminusInteger[55] = 16'b00000000_00000000;
		DminusInteger[56] = 16'b00000000_00000000;
		DminusInteger[57] = 16'b00000000_00000000;
		DminusInteger[58] = 16'b00000000_00000000;
		DminusInteger[59] = 16'b00000000_00000000;
		DminusInteger[60] = 16'b00000000_00000000;
		DminusInteger[61] = 16'b00000000_00000000;
		DminusInteger[62] = 16'b00000000_00000000;
		DminusInteger[63] = 16'b00000000_00000000;
		DminusInteger[64] = 16'b00000000_00000000;
		DminusInteger[65] = 16'b00000000_00000000;
		DminusInteger[66] = 16'b00000000_00000000;
		DminusInteger[67] = 16'b00000000_00000000;
		DminusInteger[68] = 16'b00000000_00000000;
		DminusInteger[69] = 16'b00000000_00000000;
		DminusInteger[70] = 16'b00000000_00000000;
		DminusInteger[71] = 16'b00000000_00000000;
		DminusInteger[72] = 16'b00000000_00000000;
		DminusInteger[73] = 16'b00000000_00000000;
		DminusInteger[74] = 16'b00000000_00000000;
		DminusInteger[75] = 16'b00000000_00000000;
		DminusInteger[76] = 16'b00000000_00000000;
		DminusInteger[77] = 16'b00000000_00000000;
		DminusInteger[78] = 16'b00000000_00000000;
		DminusInteger[79] = 16'b00000000_00000000;
		DminusInteger[80] = 16'b00000000_00000000;
		DminusInteger[81] = 16'b00000000_00000000;
		DminusInteger[82] = 16'b00000000_00000000;
		DminusInteger[83] = 16'b00000000_00000000;
		DminusInteger[84] = 16'b00000000_00000000;
		DminusInteger[85] = 16'b00000000_00000000;
		DminusInteger[86] = 16'b00000000_00000000;
		DminusInteger[87] = 16'b00000000_00000000;
		DminusInteger[88] = 16'b00000000_00000000;
		DminusInteger[89] = 16'b00000000_00000000;
		DminusInteger[90] = 16'b00000000_00000000;
		DminusInteger[91] = 16'b00000000_00000000;
		DminusInteger[92] = 16'b00000000_00000000;
		DminusInteger[93] = 16'b00000000_00000000;
		DminusInteger[94] = 16'b00000000_00000000;
		DminusInteger[95] = 16'b00000000_00000000;
		DminusInteger[96] = 16'b00000000_00000000;
		DminusInteger[97] = 16'b00000000_00000000;
		DminusInteger[98] = 16'b00000000_00000000;
		DminusInteger[99] = 16'b00000000_00000000;
		DminusInteger[100] = 16'b00000000_00000000;
		DminusInteger[101] = 16'b00000000_00000000;
		DminusInteger[102] = 16'b00000000_00000000;
		DminusInteger[103] = 16'b00000000_00000000;
		DminusInteger[104] = 16'b00000000_00000000;
		DminusInteger[105] = 16'b00000000_00000000;
		DminusInteger[106] = 16'b00000000_00000000;
		DminusInteger[107] = 16'b00000000_00000000;
		DminusInteger[108] = 16'b00000000_00000000;
		DminusInteger[109] = 16'b00000000_00000000;
		DminusInteger[110] = 16'b00000000_00000000;
		DminusInteger[111] = 16'b00000000_00000000;
		DminusInteger[112] = 16'b00000000_00000000;
		DminusInteger[113] = 16'b00000000_00000000;
		DminusInteger[114] = 16'b00000000_00000000;
		DminusInteger[115] = 16'b00000000_00000000;
		DminusInteger[116] = 16'b00000000_00000000;
		DminusInteger[117] = 16'b00000000_00000000;
		DminusInteger[118] = 16'b00000000_00000000;
		DminusInteger[119] = 16'b00000000_00000000;
		DminusInteger[120] = 16'b00000000_00000000;
		DminusInteger[121] = 16'b00000000_00000000;
		DminusInteger[122] = 16'b00000000_00000000;
		DminusInteger[123] = 16'b00000000_00000000;
		DminusInteger[124] = 16'b00000000_00000000;
		DminusInteger[125] = 16'b00000000_00000000;
		DminusInteger[126] = 16'b00000000_00000000;
		DminusInteger[127] = 16'b00000000_00000000;
end
endmodule
